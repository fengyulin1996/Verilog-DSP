`timescale 1ns / 1ps
module fft_top(
    input wire clk,
    input wire rstn,
    
    input wire req_i,    //fft_in
    output reg ans_o,
    input wire[15:0] data_i,
    
    input wire ans_i,    //from fft_out
    output reg req_o,
    output reg[15:0] data_oR,
    output reg[15:0] data_oJ
    );
    parameter n=10;    //点数的2的对数，即级数 n取3~10
    reg en_input,ans_input2;
    wire ans_input1_c,req_input_c;    //input_connect
    wire[15:0] data_input_c;
    
    reg en_output,req_output;
    wire req_o_c,ans_output1_c;    //output_connect
    wire[15:0] data_oR_c,data_oJ_c;
    reg[15:0] outputR,outputJ;    
    reg[15:0] a,b,c,d,e,f;
    wire[15:0] R,J;    //MAC connect
    wire over_m,over_a;
    
    reg [1:0] current_state,next_state;    //FSM
    parameter S0 = 2'b00;    //停机
    parameter S1 = 2'b01;    //输入
    parameter S2 = 2'b10;    //处理
    parameter S3 = 2'b11;    //输出
    
    
    
    reg[10:0] input_count,output_count;
    wire[10:0] vice_input_count;
    assign vice_input_count = {input_count[0],input_count[1],input_count[2],input_count[3],
                               input_count[4],input_count[5],input_count[6],input_count[7],
                               input_count[8],input_count[9]};    //码位倒序
    reg[15:0] fft0R[0:1023],fft0J[0:1023],
              fft1R[0:1023],fft1J[0:1023],fft2R[0:1023],fft2J[0:1023],
              fft3R[0:1023],fft3J[0:1023],fft4R[0:1023],fft4J[0:1023],
              fft5R[0:1023],fft5J[0:1023],fft6R[0:1023],fft6J[0:1023],
              fft7R[0:1023],fft7J[0:1023],fft8R[0:1023],fft8J[0:1023],
              fft9R[0:1023],fft9J[0:1023],fft10R[0:1023],fft10J[0:1023];
              //为蝶形运算提供运算空间，同时便于流水化
    reg[4:0] ji,next_ji;    //当前蝶形运算级（从左到右）
    reg[9:0] position,next_position,position_plus;    //当前蝶形运算位（从上到下）
    reg[15:0] W1024R[0:1023],W1024J[0:1023];    //旋转因子，在上电初始化时自动赋值
    reg[9:0] i,j;
    /*
    initial begin
    $readmemb("W1024R.dat",W1024R,0,1023);
    $readmemb("W1024J.dat",W1024J,0,1023);
    end
    */
    always @(posedge clk) begin    //状态转换
        if(rstn == 1'b0)begin
        current_state <= S0;
        
        end
        else current_state <= next_state;
    end
    always @(posedge clk) begin
        case(current_state)
            S0:begin end
            S1:begin
               fft0R[vice_input_count] <= data_input_c;
               fft0J[vice_input_count] <= 16'h0000;    //输入
               input_count = input_count + 10'b00000_00001;
               end    //S1
            S2:begin
               case(ji)
               4'b0000:begin
               
               end
               4'b0001:begin
               fft1R[position] <= R;
               fft1J[position] <= J;
               end
               4'b0010:begin
               fft2R[position] <= R;
               fft2J[position] <= J;
               end
               4'b0011:begin
               fft3R[position] <= R;
               fft3J[position] <= J;
               end
               4'b0100:begin
               fft4R[position] <= R;
               fft4J[position] <= J;
               end
               4'b0101:begin
               fft5R[position] <= R;
               fft5J[position] <= J;
               end
               4'b0110:begin
               fft6R[position] <= R;
               fft6J[position] <= J;
               end
               4'b0111:begin
               fft7R[position] <= R;
               fft7J[position] <= J;
               end
               4'b1000:begin
               fft8R[position] <= R;
               fft8J[position] <= J;
               end
               4'b1001:begin
               fft9R[position] <= R;
               fft9J[position] <= J;
               end
               4'b1010:begin
               fft10R[position] <= R;
               fft10J[position] <= J;
               end
               default:begin
               
               end
               endcase
               ji <= next_ji;    //状态转换
               position <= next_position;
               end    //S2
            S3:begin
               outputR <= fft10R[output_count];
               outputJ <= fft10J[output_count];
               output_count <= output_count + 1;
               end
        endcase
 
    end
    
    always @(*) begin    //对控制信号，次态赋值
        if(rstn == 1'b0) begin
            next_state = S0;
            input_count = 10'b00000_00000;
            
            
            
            W1024J[0] = 16'b0000000000000000;
            W1024J[1] = 16'b1111111111111110;
            W1024J[2] = 16'b1111111111111100;
            W1024J[3] = 16'b1111111111111011;
            W1024J[4] = 16'b1111111111111001;
            W1024J[5] = 16'b1111111111111000;
            W1024J[6] = 16'b1111111111110110;
            W1024J[7] = 16'b1111111111110101;
            W1024J[8] = 16'b1111111111110011;
            W1024J[9] = 16'b1111111111110001;
            W1024J[10] = 16'b1111111111110001;
            W1024J[11] = 16'b1111111111110000;
            W1024J[12] = 16'b1111111111101110;
            W1024J[13] = 16'b1111111111101101;
            W1024J[14] = 16'b1111111111101011;
            W1024J[15] = 16'b1111111111101010;
            W1024J[16] = 16'b1111111111101000;
            W1024J[17] = 16'b1111111111100110;
            W1024J[18] = 16'b1111111111100101;
            W1024J[19] = 16'b1111111111100011;
            W1024J[20] = 16'b1111111111100010;
            W1024J[21] = 16'b1111111111100000;
            W1024J[22] = 16'b1111111111011111;
            W1024J[23] = 16'b1111111111011101;
            W1024J[24] = 16'b1111111111011011;
            W1024J[25] = 16'b1111111111011010;
            W1024J[26] = 16'b1111111111011000;
            W1024J[27] = 16'b1111111111010111;
            W1024J[28] = 16'b1111111111010101;
            W1024J[29] = 16'b1111111111010100;
            W1024J[30] = 16'b1111111111010010;
            W1024J[31] = 16'b1111111111010001;
            W1024J[32] = 16'b1111111111001111;
            W1024J[33] = 16'b1111111111001110;
            W1024J[34] = 16'b1111111111001100;
            W1024J[35] = 16'b1111111111001010;
            W1024J[36] = 16'b1111111111001001;
            W1024J[37] = 16'b1111111111000111;
            W1024J[38] = 16'b1111111111000110;
            W1024J[39] = 16'b1111111111000100;
            W1024J[40] = 16'b1111111111000011;
            W1024J[41] = 16'b1111111111000001;
            W1024J[42] = 16'b1111111111000000;
            W1024J[43] = 16'b1111111110111110;
            W1024J[44] = 16'b1111111110111101;
            W1024J[45] = 16'b1111111110111011;
            W1024J[46] = 16'b1111111110111010;
            W1024J[47] = 16'b1111111110111000;
            W1024J[48] = 16'b1111111110110111;
            W1024J[49] = 16'b1111111110110101;
            W1024J[50] = 16'b1111111110110100;
            W1024J[51] = 16'b1111111110110010;
            W1024J[52] = 16'b1111111110110001;
            W1024J[53] = 16'b1111111110101111;
            W1024J[54] = 16'b1111111110101110;
            W1024J[55] = 16'b1111111110101100;
            W1024J[56] = 16'b1111111110101011;
            W1024J[57] = 16'b1111111110101001;
            W1024J[58] = 16'b1111111110101000;
            W1024J[59] = 16'b1111111110100110;
            W1024J[60] = 16'b1111111110100101;
            W1024J[61] = 16'b1111111110100011;
            W1024J[62] = 16'b1111111110100010;
            W1024J[63] = 16'b1111111110100000;
            W1024J[64] = 16'b1111111110011111;
            W1024J[65] = 16'b1111111110011110;
            W1024J[66] = 16'b1111111110011100;
            W1024J[67] = 16'b1111111110011011;
            W1024J[68] = 16'b1111111110011001;
            W1024J[69] = 16'b1111111110011000;
            W1024J[70] = 16'b1111111110010110;
            W1024J[71] = 16'b1111111110010101;
            W1024J[72] = 16'b1111111110010011;
            W1024J[73] = 16'b1111111110010010;
            W1024J[74] = 16'b1111111110010001;
            W1024J[75] = 16'b1111111110001111;
            W1024J[76] = 16'b1111111110001110;
            W1024J[77] = 16'b1111111110001100;
            W1024J[78] = 16'b1111111110001011;
            W1024J[79] = 16'b1111111110001010;
            W1024J[80] = 16'b1111111110001000;
            W1024J[81] = 16'b1111111110000111;
            W1024J[82] = 16'b1111111110000101;
            W1024J[83] = 16'b1111111110000100;
            W1024J[84] = 16'b1111111110000011;
            W1024J[85] = 16'b1111111110000001;
            W1024J[86] = 16'b1111111110000000;
            W1024J[87] = 16'b1111111101111111;
            W1024J[88] = 16'b1111111101111101;
            W1024J[89] = 16'b1111111101111100;
            W1024J[90] = 16'b1111111101111011;
            W1024J[91] = 16'b1111111101111001;
            W1024J[92] = 16'b1111111101111000;
            W1024J[93] = 16'b1111111101110111;
            W1024J[94] = 16'b1111111101110101;
            W1024J[95] = 16'b1111111101110100;
            W1024J[96] = 16'b1111111101110011;
            W1024J[97] = 16'b1111111101110001;
            W1024J[98] = 16'b1111111101110000;
            W1024J[99] = 16'b1111111101101111;
            
            W1024J[100] = 16'b1111111101101100;
            W1024J[101] = 16'b1111111101101100;
            W1024J[102] = 16'b1111111101101011;
            W1024J[103] = 16'b1111111101101010;
            W1024J[104] = 16'b1111111101101000;
            W1024J[105] = 16'b1111111101100111;
            W1024J[106] = 16'b1111111101100110;
            W1024J[107] = 16'b1111111101100100;
            W1024J[108] = 16'b1111111101100011;
            W1024J[109] = 16'b1111111101100010;
            W1024J[110] = 16'b1111111101100001;
            W1024J[111] = 16'b1111111101100000;
            W1024J[112] = 16'b1111111101011101;
            W1024J[113] = 16'b1111111101011100;
            W1024J[114] = 16'b1111111101011011;
            W1024J[115] = 16'b1111111101011001;
            W1024J[116] = 16'b1111111101011000;
            W1024J[117] = 16'b1111111101010111;
            W1024J[118] = 16'b1111111101010110;
            W1024J[119] = 16'b1111111101010101;
            W1024J[120] = 16'b1111111101010100;
            W1024J[121] = 16'b1111111101010010;
            W1024J[122] = 16'b1111111101010001;
            W1024J[123] = 16'b1111111101010000;
            W1024J[124] = 16'b1111111101001111;
            W1024J[125] = 16'b1111111101001110;
            W1024J[126] = 16'b1111111101001101;
            W1024J[127] = 16'b1111111101001100;
            W1024J[128] = 16'b1111111101001010;
            W1024J[129] = 16'b1111111101001001;
            W1024J[130] = 16'b1111111101001000;
            W1024J[131] = 16'b1111111101000111;
            W1024J[132] = 16'b1111111101000110;
            W1024J[133] = 16'b1111111101000101;
            W1024J[134] = 16'b1111111101000100;
            W1024J[135] = 16'b1111111101000011;
            W1024J[136] = 16'b1111111101000010;
            W1024J[137] = 16'b1111111101000001;
            W1024J[138] = 16'b1111111101000000;
            W1024J[139] = 16'b1111111100111111;
            W1024J[140] = 16'b1111111100111110;
            W1024J[141] = 16'b1111111100111101;
            W1024J[142] = 16'b1111111100111100;
            W1024J[143] = 16'b1111111100111011;
            W1024J[144] = 16'b1111111100111010;
            W1024J[145] = 16'b1111111100111001;
            W1024J[146] = 16'b1111111100111000;
            W1024J[147] = 16'b1111111100110111;
            W1024J[148] = 16'b1111111100110110;
            W1024J[149] = 16'b1111111100110101;
            W1024J[150] = 16'b1111111100110100;
            W1024J[151] = 16'b1111111100110011;
            W1024J[152] = 16'b1111111100110010;
            W1024J[153] = 16'b1111111100110001;
            W1024J[154] = 16'b1111111100110000;
            W1024J[155] = 16'b1111111100101111;
            W1024J[156] = 16'b1111111100101110;
            W1024J[157] = 16'b1111111100101101;
            W1024J[158] = 16'b1111111100101100;
            W1024J[159] = 16'b1111111100101100;
            W1024J[160] = 16'b1111111100101011;
            W1024J[161] = 16'b1111111100101010;
            W1024J[162] = 16'b1111111100101001;
            W1024J[163] = 16'b1111111100101000;
            W1024J[164] = 16'b1111111100100111;
            W1024J[165] = 16'b1111111100100110;
            W1024J[166] = 16'b1111111100100110;
            W1024J[167] = 16'b1111111100100101;
            W1024J[168] = 16'b1111111100100100;
            W1024J[169] = 16'b1111111100100011;
            W1024J[170] = 16'b1111111100100010;
            W1024J[171] = 16'b1111111100100010;
            W1024J[172] = 16'b1111111100100001;
            W1024J[173] = 16'b1111111100100000;
            W1024J[174] = 16'b1111111100011111;
            W1024J[175] = 16'b1111111100011110;
            W1024J[176] = 16'b1111111100011110;
            W1024J[177] = 16'b1111111100011101;
            W1024J[178] = 16'b1111111100011100;
            W1024J[179] = 16'b1111111100011100;
            W1024J[180] = 16'b1111111100011011;
            W1024J[181] = 16'b1111111100011010;
            W1024J[182] = 16'b1111111100011001;
            W1024J[183] = 16'b1111111100011001;
            W1024J[184] = 16'b1111111100011000;
            W1024J[185] = 16'b1111111100010111;
            W1024J[186] = 16'b1111111100010111;
            W1024J[187] = 16'b1111111100010110;
            W1024J[188] = 16'b1111111100010101;
            W1024J[189] = 16'b1111111100010101;
            W1024J[190] = 16'b1111111100010100;
            W1024J[191] = 16'b1111111100010100;
            W1024J[192] = 16'b1111111100010011;
            W1024J[193] = 16'b1111111100010010;
            W1024J[194] = 16'b1111111100010010;
            W1024J[195] = 16'b1111111100010010;
            W1024J[196] = 16'b1111111100010001;
            W1024J[197] = 16'b1111111100010001;
            W1024J[198] = 16'b1111111100010000;
            W1024J[199] = 16'b1111111100010000;
            
            W1024J[100+100] = 16'b1111111100001110;
            W1024J[100+101] = 16'b1111111100001110;
            W1024J[100+102] = 16'b1111111100001101;
            W1024J[100+103] = 16'b1111111100001101;
            W1024J[100+104] = 16'b1111111100001100;
            W1024J[100+105] = 16'b1111111100001100;
            W1024J[100+106] = 16'b1111111100001011;
            W1024J[100+107] = 16'b1111111100001011;
            W1024J[100+108] = 16'b1111111100001011;
            W1024J[100+109] = 16'b1111111100001010;
            W1024J[100+110] = 16'b1111111100001010;
            W1024J[100+111] = 16'b1111111100001001;
            W1024J[100+112] = 16'b1111111100001001;
            W1024J[100+113] = 16'b1111111100001000;
            W1024J[100+114] = 16'b1111111100001000;
            W1024J[100+115] = 16'b1111111100001000;
            W1024J[100+116] = 16'b1111111100000111;
            W1024J[100+117] = 16'b1111111100000111;
            W1024J[100+118] = 16'b1111111100000110;
            W1024J[100+119] = 16'b1111111100000110;
            W1024J[100+120] = 16'b1111111100000110;
            W1024J[100+121] = 16'b1111111100000101;
            W1024J[100+122] = 16'b1111111100000101;
            W1024J[100+123] = 16'b1111111100000101;
            W1024J[100+124] = 16'b1111111100000100;
            W1024J[100+125] = 16'b1111111100000100;
            W1024J[100+126] = 16'b1111111100000100;
            W1024J[100+127] = 16'b1111111100000100;
            W1024J[100+128] = 16'b1111111100000011;
            W1024J[100+129] = 16'b1111111100000011;
            W1024J[100+130] = 16'b1111111100000011;
            W1024J[100+131] = 16'b1111111100000011;
            W1024J[100+132] = 16'b1111111100000010;
            W1024J[100+133] = 16'b1111111100000010;
            W1024J[100+134] = 16'b1111111100000010;
            W1024J[100+135] = 16'b1111111100000010;
            W1024J[100+136] = 16'b1111111100000001;
            W1024J[100+137] = 16'b1111111100000001;
            W1024J[100+138] = 16'b1111111100000001;
            W1024J[100+139] = 16'b1111111100000001;
            W1024J[100+140] = 16'b1111111100000001;
            W1024J[100+141] = 16'b1111111100000001;
            W1024J[100+142] = 16'b1111111100000001;
            W1024J[100+143] = 16'b1111111100000000;
            W1024J[100+144] = 16'b1111111100000000;
            W1024J[100+145] = 16'b1111111100000000;
            W1024J[100+146] = 16'b1111111100000000;
            W1024J[100+147] = 16'b1111111100000000;
            W1024J[100+148] = 16'b1111111100000000;
            W1024J[100+149] = 16'b1111111100000000;
            W1024J[100+150] = 16'b1111111100000000;
            W1024J[100+151] = 16'b1111111100000000;
            W1024J[100+152] = 16'b1111111100000000;
            W1024J[100+153] = 16'b1111111100000000;
            W1024J[100+154] = 16'b1111111100000000;
            W1024J[100+155] = 16'b1111111100000000;
            W1024J[100+156] = 16'b1111111100000000;
            W1024J[100+157] = 16'b1111111100000000;
            W1024J[100+158] = 16'b1111111100000000;
            W1024J[100+159] = 16'b1111111100000000;
            W1024J[100+160] = 16'b1111111100000000;
            W1024J[100+161] = 16'b1111111100000000;
            W1024J[100+162] = 16'b1111111100000000;
            W1024J[100+163] = 16'b1111111100000000;
            W1024J[100+164] = 16'b1111111100000000;
            W1024J[100+165] = 16'b1111111100000000;
            W1024J[100+166] = 16'b1111111100000000;
            W1024J[100+167] = 16'b1111111100000000;
            W1024J[100+168] = 16'b1111111100000000;
            W1024J[100+169] = 16'b1111111100000000;
            W1024J[100+170] = 16'b1111111100000000;
            W1024J[100+171] = 16'b1111111100000000;
            W1024J[100+172] = 16'b1111111100000001;
            W1024J[100+173] = 16'b1111111100000001;
            W1024J[100+174] = 16'b1111111100000001;
            W1024J[100+175] = 16'b1111111100000001;
            W1024J[100+176] = 16'b1111111100000001;
            W1024J[100+177] = 16'b1111111100000001;
            W1024J[100+178] = 16'b1111111100000010;
            W1024J[100+179] = 16'b1111111100000010;
            W1024J[100+180] = 16'b1111111100000010;
            W1024J[100+181] = 16'b1111111100000010;
            W1024J[100+182] = 16'b1111111100000011;
            W1024J[100+183] = 16'b1111111100000011;
            W1024J[100+184] = 16'b1111111100000011;
            W1024J[100+185] = 16'b1111111100000011;
            W1024J[100+186] = 16'b1111111100000100;
            W1024J[100+187] = 16'b1111111100000100;
            W1024J[100+188] = 16'b1111111100000100;
            W1024J[100+189] = 16'b1111111100000100;
            W1024J[100+190] = 16'b1111111100000101;
            W1024J[100+191] = 16'b1111111100000101;
            W1024J[100+192] = 16'b1111111100000101;
            W1024J[100+193] = 16'b1111111100000110;
            W1024J[100+194] = 16'b1111111100000110;
            W1024J[100+195] = 16'b1111111100000110;
            W1024J[100+196] = 16'b1111111100000111;
            W1024J[100+197] = 16'b1111111100000111;
            W1024J[100+198] = 16'b1111111100001000;
            W1024J[100+199] = 16'b1111111100001000;
            
            
            
            W1024J[200+100] = 16'b1111111100001001;
            W1024J[200+101] = 16'b1111111100001001;
            W1024J[200+102] = 16'b1111111100001010;
            W1024J[200+103] = 16'b1111111100001010;
            W1024J[200+104] = 16'b1111111100001011;
            W1024J[200+105] = 16'b1111111100001011;
            W1024J[200+106] = 16'b1111111100001011;
            W1024J[200+107] = 16'b1111111100001100;
            W1024J[200+108] = 16'b1111111100001100;
            W1024J[200+109] = 16'b1111111100001101;
            W1024J[200+110] = 16'b1111111100001101;
            W1024J[200+111] = 16'b1111111100001110;
            W1024J[200+112] = 16'b1111111100001110;
            W1024J[200+113] = 16'b1111111100001111;
            W1024J[200+114] = 16'b1111111100010000;
            W1024J[200+115] = 16'b1111111100010000;
            W1024J[200+116] = 16'b1111111100010001;
            W1024J[200+117] = 16'b1111111100010001;
            W1024J[200+118] = 16'b1111111100010010;
            W1024J[200+119] = 16'b1111111100010010;
            W1024J[200+120] = 16'b1111111100010011;
            W1024J[200+121] = 16'b1111111100010100;
            W1024J[200+122] = 16'b1111111100010100;
            W1024J[200+123] = 16'b1111111100010101;
            W1024J[200+124] = 16'b1111111100010101;
            W1024J[200+125] = 16'b1111111100010110;
            W1024J[200+126] = 16'b1111111100010111;
            W1024J[200+127] = 16'b1111111100010111;
            W1024J[200+128] = 16'b1111111100011000;
            W1024J[200+129] = 16'b1111111100011001;
            W1024J[200+130] = 16'b1111111100011001;
            W1024J[200+131] = 16'b1111111100011010;
            W1024J[200+132] = 16'b1111111100011011;
            W1024J[200+133] = 16'b1111111100011100;
            W1024J[200+134] = 16'b1111111100011100;
            W1024J[200+135] = 16'b1111111100011101;
            W1024J[200+136] = 16'b1111111100011110;
            W1024J[200+137] = 16'b1111111100011110;
            W1024J[200+138] = 16'b1111111100011111;
            W1024J[200+139] = 16'b1111111100100000;
            W1024J[200+140] = 16'b1111111100100001;
            W1024J[200+141] = 16'b1111111100100010;
            W1024J[200+142] = 16'b1111111100100010;
            W1024J[200+143] = 16'b1111111100100011;
            W1024J[200+144] = 16'b1111111100100100;
            W1024J[200+145] = 16'b1111111100100101;
            W1024J[200+146] = 16'b1111111100100110;
            W1024J[200+147] = 16'b1111111100100110;
            W1024J[200+148] = 16'b1111111100100111;
            W1024J[200+149] = 16'b1111111100100110;
            W1024J[200+150] = 16'b1111111100100111;
            W1024J[200+151] = 16'b1111111100101000;
            W1024J[200+152] = 16'b1111111100101001;
            W1024J[200+153] = 16'b1111111100101010;
            W1024J[200+154] = 16'b1111111100101011;
            W1024J[200+155] = 16'b1111111100101100;
            W1024J[200+156] = 16'b1111111100101100;
            W1024J[200+157] = 16'b1111111100101101;
            W1024J[200+158] = 16'b1111111100101110;
            W1024J[200+159] = 16'b1111111100101111;
            W1024J[200+160] = 16'b1111111100110000;
            W1024J[200+161] = 16'b1111111100110001;
            W1024J[200+162] = 16'b1111111100110010;
            W1024J[200+163] = 16'b1111111100110011;
            W1024J[200+164] = 16'b1111111100110100;
            W1024J[200+165] = 16'b1111111100110101;
            W1024J[200+166] = 16'b1111111100110111;
            W1024J[200+167] = 16'b1111111100111000;
            W1024J[200+168] = 16'b1111111100111001;
            W1024J[200+169] = 16'b1111111100111010;
            W1024J[200+170] = 16'b1111111100111011;
            W1024J[200+171] = 16'b1111111100111100;
            W1024J[200+172] = 16'b1111111100111101;
            W1024J[200+173] = 16'b1111111100111110;
            W1024J[200+174] = 16'b1111111100111111;
            W1024J[200+175] = 16'b1111111101000000;
            W1024J[200+176] = 16'b1111111101000001;
            W1024J[200+177] = 16'b1111111101000010;
            W1024J[200+178] = 16'b1111111101000011;
            W1024J[200+179] = 16'b1111111101000100;
            W1024J[200+180] = 16'b1111111101000101;
            W1024J[200+181] = 16'b1111111101000110;
            W1024J[200+182] = 16'b1111111101000111;
            W1024J[200+183] = 16'b1111111101001000;
            W1024J[200+184] = 16'b1111111101001001;
            W1024J[200+185] = 16'b1111111101001010;
            W1024J[200+186] = 16'b1111111101001100;
            W1024J[200+187] = 16'b1111111101001101;
            W1024J[200+188] = 16'b1111111101001110;
            W1024J[200+189] = 16'b1111111101001111;
            W1024J[200+190] = 16'b1111111101010000;
            W1024J[200+191] = 16'b1111111101010001;
            W1024J[200+192] = 16'b1111111101010010;
            W1024J[200+193] = 16'b1111111101010100;
            W1024J[200+194] = 16'b1111111101010101;
            W1024J[200+195] = 16'b1111111101010110;
            W1024J[200+196] = 16'b1111111101010111;
            W1024J[200+197] = 16'b1111111101011000;
            W1024J[200+198] = 16'b1111111101011001;
            W1024J[200+199] = 16'b1111111101011011;
            
            W1024J[300+100] = 16'b0000_0001_0000_0000;
            W1024J[300+101] = 16'b0000_0001_0000_0000;
            W1024J[300+102] = 16'b0000_0001_0000_0000;
            W1024J[300+103] = 16'b0000_0001_0000_0000;
            W1024J[300+104] = 16'b0000_0001_0000_0000;
            W1024J[300+105] = 16'b0000_0001_0000_0000;
            W1024J[300+106] = 16'b0000_0001_0000_0000;
            W1024J[300+107] = 16'b0000_0001_0000_0000;
            W1024J[300+108] = 16'b0000_0001_0000_0000;
            W1024J[300+109] = 16'b0000_0001_0000_0000;
            W1024J[300+110] = 16'b0000_0001_0000_0000;
            W1024J[300+111] = 16'b0000_0001_0000_0000;
            W1024J[300+112] = 16'b0000_0001_0000_0000;
            W1024J[300+113] = 16'b0000_0001_0000_0000;
            W1024J[300+114] = 16'b0000_0001_0000_0000;
            W1024J[300+115] = 16'b0000_0001_0000_0000;
            W1024J[300+116] = 16'b0000_0001_0000_0000;
            W1024J[300+117] = 16'b0000_0001_0000_0000;
            W1024J[300+118] = 16'b0000_0001_0000_0000;
            W1024J[300+119] = 16'b0000_0001_0000_0000;
            W1024J[300+120] = 16'b0000_0001_0000_0000;
            W1024J[300+121] = 16'b0000_0001_0000_0000;
            W1024J[300+122] = 16'b0000_0001_0000_0000;
            W1024J[300+123] = 16'b0000_0001_0000_0000;
            W1024J[300+124] = 16'b0000_0001_0000_0000;
            W1024J[300+125] = 16'b0000_0001_0000_0000;
            W1024J[300+126] = 16'b0000_0001_0000_0000;
            W1024J[300+127] = 16'b0000_0001_0000_0000;
            W1024J[300+128] = 16'b0000_0001_0000_0000;
            W1024J[300+129] = 16'b0000_0001_0000_0000;
            W1024J[300+130] = 16'b0000_0001_0000_0000;
            W1024J[300+131] = 16'b0000_0001_0000_0000;
            W1024J[300+132] = 16'b0000_0001_0000_0000;
            W1024J[300+133] = 16'b0000_0001_0000_0000;
            W1024J[300+134] = 16'b0000_0001_0000_0000;
            W1024J[300+135] = 16'b0000_0001_0000_0000;
            W1024J[300+136] = 16'b0000_0001_0000_0000;
            W1024J[300+137] = 16'b0000_0001_0000_0000;
            W1024J[300+138] = 16'b0000_0001_0000_0000;
            W1024J[300+139] = 16'b0000_0001_0000_0000;
            W1024J[300+140] = 16'b0000_0001_0000_0000;
            W1024J[300+141] = 16'b0000_0001_0000_0000;
            W1024J[300+142] = 16'b0000_0001_0000_0000;
            W1024J[300+143] = 16'b0000_0001_0000_0000;
            W1024J[300+144] = 16'b0000_0001_0000_0000;
            W1024J[300+145] = 16'b0000_0001_0000_0000;
            W1024J[300+146] = 16'b0000_0001_0000_0000;
            W1024J[300+147] = 16'b0000_0001_0000_0000;
            W1024J[300+148] = 16'b0000_0001_0000_0000;
            W1024J[300+149] = 16'b0000_0001_0000_0000;
            W1024J[300+150] = 16'b0000_0001_0000_0000;
            W1024J[300+151] = 16'b0000_0001_0000_0000;
            W1024J[300+152] = 16'b0000_0001_0000_0000;
            W1024J[300+153] = 16'b0000_0001_0000_0000;
            W1024J[300+154] = 16'b0000_0001_0000_0000;
            W1024J[300+155] = 16'b0000_0001_0000_0000;
            W1024J[300+156] = 16'b0000_0001_0000_0000;
            W1024J[300+157] = 16'b0000_0001_0000_0000;
            W1024J[300+158] = 16'b0000_0001_0000_0000;
            W1024J[300+159] = 16'b0000_0001_0000_0000;
            W1024J[300+160] = 16'b0000_0001_0000_0000;
            W1024J[300+161] = 16'b0000_0001_0000_0000;
            W1024J[300+162] = 16'b0000_0001_0000_0000;
            W1024J[300+163] = 16'b0000_0001_0000_0000;
            W1024J[300+164] = 16'b0000_0001_0000_0000;
            W1024J[300+165] = 16'b0000_0001_0000_0000;
            W1024J[300+166] = 16'b0000_0001_0000_0000;
            W1024J[300+167] = 16'b0000_0001_0000_0000;
            W1024J[300+168] = 16'b0000_0001_0000_0000;
            W1024J[300+169] = 16'b0000_0001_0000_0000;
            W1024J[300+170] = 16'b0000_0001_0000_0000;
            W1024J[300+171] = 16'b0000_0001_0000_0000;
            W1024J[300+172] = 16'b0000_0001_0000_0000;
            W1024J[300+173] = 16'b0000_0001_0000_0000;
            W1024J[300+174] = 16'b0000_0001_0000_0000;
            W1024J[300+175] = 16'b0000_0001_0000_0000;
            W1024J[300+176] = 16'b0000_0001_0000_0000;
            W1024J[300+177] = 16'b0000_0001_0000_0000;
            W1024J[300+178] = 16'b0000_0001_0000_0000;
            W1024J[300+179] = 16'b0000_0001_0000_0000;
            W1024J[300+180] = 16'b0000_0001_0000_0000;
            W1024J[300+181] = 16'b0000_0001_0000_0000;
            W1024J[300+182] = 16'b0000_0001_0000_0000;
            W1024J[300+183] = 16'b0000_0001_0000_0000;
            W1024J[300+184] = 16'b0000_0001_0000_0000;
            W1024J[300+185] = 16'b0000_0001_0000_0000;
            W1024J[300+186] = 16'b0000_0001_0000_0000;
            W1024J[300+187] = 16'b0000_0001_0000_0000;
            W1024J[300+188] = 16'b0000_0001_0000_0000;
            W1024J[300+189] = 16'b0000_0001_0000_0000;
            W1024J[300+190] = 16'b0000_0001_0000_0000;
            W1024J[300+191] = 16'b0000_0001_0000_0000;
            W1024J[300+192] = 16'b0000_0001_0000_0000;
            W1024J[300+193] = 16'b0000_0001_0000_0000;
            W1024J[300+194] = 16'b0000_0001_0000_0000;
            W1024J[300+195] = 16'b0000_0001_0000_0000;
            W1024J[300+196] = 16'b0000_0001_0000_0000;
            W1024J[300+197] = 16'b0000_0001_0000_0000;
            W1024J[300+198] = 16'b0000_0001_0000_0000;
            W1024J[300+199] = 16'b0000_0001_0000_0000;
            
            W1024J[400+100] = 16'b0000_0001_0000_0000;
            W1024J[400+101] = 16'b0000_0001_0000_0000;
            W1024J[400+102] = 16'b0000_0001_0000_0000;
            W1024J[400+103] = 16'b0000_0001_0000_0000;
            W1024J[400+104] = 16'b0000_0001_0000_0000;
            W1024J[400+105] = 16'b0000_0001_0000_0000;
            W1024J[400+106] = 16'b0000_0001_0000_0000;
            W1024J[400+107] = 16'b0000_0001_0000_0000;
            W1024J[400+108] = 16'b0000_0001_0000_0000;
            W1024J[400+109] = 16'b0000_0001_0000_0000;
            W1024J[400+110] = 16'b0000_0001_0000_0000;
            W1024J[400+111] = 16'b0000_0001_0000_0000;
            W1024J[400+112] = 16'b0000_0001_0000_0000;
            
            

            W1024J[400+113] = 16'b0000_0001_0000_0000;
            W1024J[400+114] = 16'b0000_0001_0000_0000;
            W1024J[400+115] = 16'b0000_0001_0000_0000;
            W1024J[400+116] = 16'b0000_0001_0000_0000;
            W1024J[400+117] = 16'b0000_0001_0000_0000;
            W1024J[400+118] = 16'b0000_0001_0000_0000;
            W1024J[400+119] = 16'b0000_0001_0000_0000;
            W1024J[400+120] = 16'b0000_0001_0000_0000;
            W1024J[400+121] = 16'b0000_0001_0000_0000;
            W1024J[400+122] = 16'b0000_0001_0000_0000;
            W1024J[400+123] = 16'b0000_0001_0000_0000;
            W1024J[400+124] = 16'b0000_0001_0000_0000;
            W1024J[400+125] = 16'b0000_0001_0000_0000;
            W1024J[400+126] = 16'b0000_0001_0000_0000;
            W1024J[400+127] = 16'b0000_0001_0000_0000;
            W1024J[400+128] = 16'b0000_0001_0000_0000;
            W1024J[400+129] = 16'b0000_0001_0000_0000;
            W1024J[400+130] = 16'b0000_0001_0000_0000;
            W1024J[400+131] = 16'b0000_0001_0000_0000;
            W1024J[400+132] = 16'b0000_0001_0000_0000;
            W1024J[400+133] = 16'b0000_0001_0000_0000;
            W1024J[400+134] = 16'b0000_0001_0000_0000;
            W1024J[400+135] = 16'b0000_0001_0000_0000;
            W1024J[400+136] = 16'b0000_0001_0000_0000;
            W1024J[400+137] = 16'b0000_0001_0000_0000;
            W1024J[400+138] = 16'b0000_0001_0000_0000;
            W1024J[400+139] = 16'b0000_0001_0000_0000;
            W1024J[400+140] = 16'b0000_0001_0000_0000;
            W1024J[400+141] = 16'b0000_0001_0000_0000;
            W1024J[400+142] = 16'b0000_0001_0000_0000;
            W1024J[400+143] = 16'b0000_0001_0000_0000;
            W1024J[400+144] = 16'b0000_0001_0000_0000;
            W1024J[400+145] = 16'b0000_0001_0000_0000;
            W1024J[400+146] = 16'b0000_0001_0000_0000;
            W1024J[400+147] = 16'b0000_0001_0000_0000;
            W1024J[400+148] = 16'b0000_0001_0000_0000;
            W1024J[400+149] = 16'b0000_0001_0000_0000;
            W1024J[400+150] = 16'b0000_0001_0000_0000;
            W1024J[400+151] = 16'b0000_0001_0000_0000;
            W1024J[400+152] = 16'b0000_0001_0000_0000;
            W1024J[400+153] = 16'b0000_0001_0000_0000;
            W1024J[400+154] = 16'b0000_0001_0000_0000;
            W1024J[400+155] = 16'b0000_0001_0000_0000;
            W1024J[400+156] = 16'b0000_0001_0000_0000;
            W1024J[400+157] = 16'b0000_0001_0000_0000;
            W1024J[400+158] = 16'b0000_0001_0000_0000;
            W1024J[400+159] = 16'b0000_0001_0000_0000;
            W1024J[400+160] = 16'b0000_0001_0000_0000;
            W1024J[400+161] = 16'b0000_0001_0000_0000;
            W1024J[400+162] = 16'b0000_0001_0000_0000;
            W1024J[400+163] = 16'b0000_0001_0000_0000;
            W1024J[400+164] = 16'b0000_0001_0000_0000;
            W1024J[400+165] = 16'b0000_0001_0000_0000;
            W1024J[400+166] = 16'b0000_0001_0000_0000;
            W1024J[400+167] = 16'b0000_0001_0000_0000;
            W1024J[400+168] = 16'b0000_0001_0000_0000;
            W1024J[400+169] = 16'b0000_0001_0000_0000;
            W1024J[400+170] = 16'b0000_0001_0000_0000;
            W1024J[400+171] = 16'b0000_0001_0000_0000;
            W1024J[400+172] = 16'b0000_0001_0000_0000;
            W1024J[400+173] = 16'b0000_0001_0000_0000;
            W1024J[400+174] = 16'b0000_0001_0000_0000;
            W1024J[400+175] = 16'b0000_0001_0000_0000;
            W1024J[400+176] = 16'b0000_0001_0000_0000;
            W1024J[400+177] = 16'b0000_0001_0000_0000;
            W1024J[400+178] = 16'b0000_0001_0000_0000;
            W1024J[400+179] = 16'b0000_0001_0000_0000;
            W1024J[400+180] = 16'b0000_0001_0000_0000;
            W1024J[400+181] = 16'b0000_0001_0000_0000;
            W1024J[400+182] = 16'b0000_0001_0000_0000;
            W1024J[400+183] = 16'b0000_0001_0000_0000;
            W1024J[400+184] = 16'b0000_0001_0000_0000;
            W1024J[400+185] = 16'b0000_0001_0000_0000;
            W1024J[400+186] = 16'b0000_0001_0000_0000;
            W1024J[400+187] = 16'b0000_0001_0000_0000;
            W1024J[400+188] = 16'b0000_0001_0000_0000;
            W1024J[400+189] = 16'b0000_0001_0000_0000;
            W1024J[400+190] = 16'b0000_0001_0000_0000;
            W1024J[400+191] = 16'b0000_0001_0000_0000;
            W1024J[400+192] = 16'b0000_0001_0000_0000;
            W1024J[400+193] = 16'b0000_0001_0000_0000;
            W1024J[400+194] = 16'b0000_0001_0000_0000;
            W1024J[400+195] = 16'b0000_0001_0000_0000;
            W1024J[400+196] = 16'b0000_0001_0000_0000;
            W1024J[400+197] = 16'b0000_0001_0000_0000;
            W1024J[400+198] = 16'b0000_0001_0000_0000;
            W1024J[400+199] = 16'b0000_0001_0000_0000;
            
            W1024J[500+100] = 16'b0000_0001_0000_0000;
            W1024J[500+101] = 16'b0000_0001_0000_0000;
            W1024J[500+102] = 16'b0000_0001_0000_0000;
            W1024J[500+103] = 16'b0000_0001_0000_0000;
            W1024J[500+104] = 16'b0000_0001_0000_0000;
            W1024J[500+105] = 16'b0000_0001_0000_0000;
            W1024J[500+106] = 16'b0000_0001_0000_0000;
            W1024J[500+107] = 16'b0000_0001_0000_0000;
            W1024J[500+108] = 16'b0000_0001_0000_0000;
            W1024J[500+109] = 16'b0000_0001_0000_0000;
            W1024J[500+110] = 16'b0000_0001_0000_0000;
            W1024J[500+111] = 16'b0000_0001_0000_0000;
            W1024J[500+112] = 16'b0000_0001_0000_0000;
            W1024J[500+113] = 16'b0000_0001_0000_0000;
            W1024J[500+114] = 16'b0000_0001_0000_0000;
            W1024J[500+115] = 16'b0000_0001_0000_0000;
            W1024J[500+116] = 16'b0000_0001_0000_0000;
            W1024J[500+117] = 16'b0000_0001_0000_0000;
            W1024J[500+118] = 16'b0000_0001_0000_0000;
            W1024J[500+119] = 16'b0000_0001_0000_0000;
            W1024J[500+120] = 16'b0000_0001_0000_0000;
            W1024J[500+121] = 16'b0000_0001_0000_0000;
            W1024J[500+122] = 16'b0000_0001_0000_0000;
            W1024J[500+123] = 16'b0000_0001_0000_0000;
            W1024J[500+124] = 16'b0000_0001_0000_0000;
            W1024J[500+125] = 16'b0000_0001_0000_0000;
            W1024J[500+126] = 16'b0000_0001_0000_0000;
            W1024J[500+127] = 16'b0000_0001_0000_0000;
            W1024J[500+128] = 16'b0000_0001_0000_0000;
            W1024J[500+129] = 16'b0000_0001_0000_0000;
            W1024J[500+130] = 16'b0000_0001_0000_0000;
            W1024J[500+131] = 16'b0000_0001_0000_0000;
            W1024J[500+132] = 16'b0000_0001_0000_0000;
            W1024J[500+133] = 16'b0000_0001_0000_0000;
            W1024J[500+134] = 16'b0000_0001_0000_0000;
            W1024J[500+135] = 16'b0000_0001_0000_0000;
            W1024J[500+136] = 16'b0000_0001_0000_0000;
            W1024J[500+137] = 16'b0000_0001_0000_0000;
            W1024J[500+138] = 16'b0000_0001_0000_0000;
            W1024J[500+139] = 16'b0000_0001_0000_0000;
            W1024J[500+140] = 16'b0000_0001_0000_0000;
            W1024J[500+141] = 16'b0000_0001_0000_0000;
            W1024J[500+142] = 16'b0000_0001_0000_0000;
            W1024J[500+143] = 16'b0000_0001_0000_0000;
            W1024J[500+144] = 16'b0000_0001_0000_0000;
            W1024J[500+145] = 16'b0000_0001_0000_0000;
            W1024J[500+146] = 16'b0000_0001_0000_0000;
            W1024J[500+147] = 16'b0000_0001_0000_0000;
            W1024J[500+148] = 16'b0000_0001_0000_0000;
            W1024J[500+149] = 16'b0000_0001_0000_0000;
            W1024J[500+150] = 16'b0000_0001_0000_0000;
            W1024J[500+151] = 16'b0000_0001_0000_0000;
            W1024J[500+152] = 16'b0000_0001_0000_0000;
            W1024J[500+153] = 16'b0000_0001_0000_0000;
            W1024J[500+154] = 16'b0000_0001_0000_0000;
            W1024J[500+155] = 16'b0000_0001_0000_0000;
            W1024J[500+156] = 16'b0000_0001_0000_0000;
            W1024J[500+157] = 16'b0000_0001_0000_0000;
            W1024J[500+158] = 16'b0000_0001_0000_0000;
            W1024J[500+159] = 16'b0000_0001_0000_0000;
            W1024J[500+160] = 16'b0000_0001_0000_0000;
            W1024J[500+161] = 16'b0000_0001_0000_0000;
            W1024J[500+162] = 16'b0000_0001_0000_0000;
            W1024J[500+163] = 16'b0000_0001_0000_0000;
            W1024J[500+164] = 16'b0000_0001_0000_0000;
            W1024J[500+165] = 16'b0000_0001_0000_0000;
            W1024J[500+166] = 16'b0000_0001_0000_0000;
            W1024J[500+167] = 16'b0000_0001_0000_0000;
            W1024J[500+168] = 16'b0000_0001_0000_0000;
            W1024J[500+169] = 16'b0000_0001_0000_0000;
            W1024J[500+170] = 16'b0000_0001_0000_0000;
            W1024J[500+171] = 16'b0000_0001_0000_0000;
            W1024J[500+172] = 16'b0000_0001_0000_0000;
            W1024J[500+173] = 16'b0000_0001_0000_0000;
            W1024J[500+174] = 16'b0000_0001_0000_0000;
            W1024J[500+175] = 16'b0000_0001_0000_0000;
            W1024J[500+176] = 16'b0000_0001_0000_0000;
            W1024J[500+177] = 16'b0000_0001_0000_0000;
            W1024J[500+178] = 16'b0000_0001_0000_0000;
            W1024J[500+179] = 16'b0000_0001_0000_0000;
            W1024J[500+180] = 16'b0000_0001_0000_0000;
            W1024J[500+181] = 16'b0000_0001_0000_0000;
            W1024J[500+182] = 16'b0000_0001_0000_0000;
            W1024J[500+183] = 16'b0000_0001_0000_0000;
            W1024J[500+184] = 16'b0000_0001_0000_0000;
            W1024J[500+185] = 16'b0000_0001_0000_0000;
            W1024J[500+186] = 16'b0000_0001_0000_0000;
            W1024J[500+187] = 16'b0000_0001_0000_0000;
            W1024J[500+188] = 16'b0000_0001_0000_0000;
            W1024J[500+189] = 16'b0000_0001_0000_0000;
            W1024J[500+190] = 16'b0000_0001_0000_0000;
            W1024J[500+191] = 16'b0000_0001_0000_0000;
            W1024J[500+192] = 16'b0000_0001_0000_0000;
            W1024J[500+193] = 16'b0000_0001_0000_0000;
            W1024J[500+194] = 16'b0000_0001_0000_0000;
            W1024J[500+195] = 16'b0000_0001_0000_0000;
            W1024J[500+196] = 16'b0000_0001_0000_0000;
            W1024J[500+197] = 16'b0000_0001_0000_0000;
            W1024J[500+198] = 16'b0000_0001_0000_0000;
            W1024J[500+199] = 16'b0000_0001_0000_0000;
            
            W1024J[600+100] = 16'b0000_0001_0000_0000;
            W1024J[600+101] = 16'b0000_0001_0000_0000;
            W1024J[600+102] = 16'b0000_0001_0000_0000;
            W1024J[600+103] = 16'b0000_0001_0000_0000;
            W1024J[600+104] = 16'b0000_0001_0000_0000;
            W1024J[600+105] = 16'b0000_0001_0000_0000;
            W1024J[600+106] = 16'b0000_0001_0000_0000;
            W1024J[600+107] = 16'b0000_0001_0000_0000;
            W1024J[600+108] = 16'b0000_0001_0000_0000;
            W1024J[600+109] = 16'b0000_0001_0000_0000;
            W1024J[600+110] = 16'b0000_0001_0000_0000;
            W1024J[600+111] = 16'b0000_0001_0000_0000;
            W1024J[600+112] = 16'b0000_0001_0000_0000;
            W1024J[600+113] = 16'b0000_0001_0000_0000;
            W1024J[600+114] = 16'b0000_0001_0000_0000;
            W1024J[600+115] = 16'b0000_0001_0000_0000;
            W1024J[600+116] = 16'b0000_0001_0000_0000;
            W1024J[600+117] = 16'b0000_0001_0000_0000;
            W1024J[600+118] = 16'b0000_0001_0000_0000;
            W1024J[600+119] = 16'b0000_0001_0000_0000;
            W1024J[600+120] = 16'b0000_0001_0000_0000;
            W1024J[600+121] = 16'b0000_0001_0000_0000;
            W1024J[600+122] = 16'b0000_0001_0000_0000;
            W1024J[600+123] = 16'b0000_0001_0000_0000;
            W1024J[600+124] = 16'b0000_0001_0000_0000;
            W1024J[600+125] = 16'b0000_0001_0000_0000;
            W1024J[600+126] = 16'b0000_0001_0000_0000;
            W1024J[600+127] = 16'b0000_0001_0000_0000;
            W1024J[600+128] = 16'b0000_0001_0000_0000;
            W1024J[600+129] = 16'b0000_0001_0000_0000;
            W1024J[600+130] = 16'b0000_0001_0000_0000;
            W1024J[600+131] = 16'b0000_0001_0000_0000;
            W1024J[600+132] = 16'b0000_0001_0000_0000;
            W1024J[600+133] = 16'b0000_0001_0000_0000;
            W1024J[600+134] = 16'b0000_0001_0000_0000;
            W1024J[600+135] = 16'b0000_0001_0000_0000;
            W1024J[600+136] = 16'b0000_0001_0000_0000;
            W1024J[600+137] = 16'b0000_0001_0000_0000;
            W1024J[600+138] = 16'b0000_0001_0000_0000;
            W1024J[600+139] = 16'b0000_0001_0000_0000;
            W1024J[600+140] = 16'b0000_0001_0000_0000;
            W1024J[600+141] = 16'b0000_0001_0000_0000;
            W1024J[600+142] = 16'b0000_0001_0000_0000;
            W1024J[600+143] = 16'b0000_0001_0000_0000;
            W1024J[600+144] = 16'b0000_0001_0000_0000;
            W1024J[600+145] = 16'b0000_0001_0000_0000;
            W1024J[600+146] = 16'b0000_0001_0000_0000;
            W1024J[600+147] = 16'b0000_0001_0000_0000;
            W1024J[600+148] = 16'b0000_0001_0000_0000;
            W1024J[600+149] = 16'b0000_0001_0000_0000;
            W1024J[600+150] = 16'b0000_0001_0000_0000;
            W1024J[600+151] = 16'b0000_0001_0000_0000;
            W1024J[600+152] = 16'b0000_0001_0000_0000;
            W1024J[600+153] = 16'b0000_0001_0000_0000;
            W1024J[600+154] = 16'b0000_0001_0000_0000;
            W1024J[600+155] = 16'b0000_0001_0000_0000;
            W1024J[600+156] = 16'b0000_0001_0000_0000;
            W1024J[600+157] = 16'b0000_0001_0000_0000;
            W1024J[600+158] = 16'b0000_0001_0000_0000;
            W1024J[600+159] = 16'b0000_0001_0000_0000;
            W1024J[600+160] = 16'b0000_0001_0000_0000;
            W1024J[600+161] = 16'b0000_0001_0000_0000;
            W1024J[600+162] = 16'b0000_0001_0000_0000;
            W1024J[600+163] = 16'b0000_0001_0000_0000;
            W1024J[600+164] = 16'b0000_0001_0000_0000;
            W1024J[600+165] = 16'b0000_0001_0000_0000;
            W1024J[600+166] = 16'b0000_0001_0000_0000;
            W1024J[600+167] = 16'b0000_0001_0000_0000;
            W1024J[600+168] = 16'b0000_0001_0000_0000;
            W1024J[600+169] = 16'b0000_0001_0000_0000;
            W1024J[600+170] = 16'b0000_0001_0000_0000;
            W1024J[600+171] = 16'b0000_0001_0000_0000;
            W1024J[600+172] = 16'b0000_0001_0000_0000;
            W1024J[600+173] = 16'b0000_0001_0000_0000;
            W1024J[600+174] = 16'b0000_0001_0000_0000;
            W1024J[600+175] = 16'b0000_0001_0000_0000;
            W1024J[600+176] = 16'b0000_0001_0000_0000;
            W1024J[600+177] = 16'b0000_0001_0000_0000;
            W1024J[600+178] = 16'b0000_0001_0000_0000;
            W1024J[600+179] = 16'b0000_0001_0000_0000;
            W1024J[600+180] = 16'b0000_0001_0000_0000;
            W1024J[600+181] = 16'b0000_0001_0000_0000;
            W1024J[600+182] = 16'b0000_0001_0000_0000;
            W1024J[600+183] = 16'b0000_0001_0000_0000;
            W1024J[600+184] = 16'b0000_0001_0000_0000;
            W1024J[600+185] = 16'b0000_0001_0000_0000;
            W1024J[600+186] = 16'b0000_0001_0000_0000;
            W1024J[600+187] = 16'b0000_0001_0000_0000;
            W1024J[600+188] = 16'b0000_0001_0000_0000;
            W1024J[600+189] = 16'b0000_0001_0000_0000;
            W1024J[600+190] = 16'b0000_0001_0000_0000;
            W1024J[600+191] = 16'b0000_0001_0000_0000;
            W1024J[600+192] = 16'b0000_0001_0000_0000;
            W1024J[600+193] = 16'b0000_0001_0000_0000;
            W1024J[600+194] = 16'b0000_0001_0000_0000;
            W1024J[600+195] = 16'b0000_0001_0000_0000;
            W1024J[600+196] = 16'b0000_0001_0000_0000;
            W1024J[600+197] = 16'b0000_0001_0000_0000;
            W1024J[600+198] = 16'b0000_0001_0000_0000;
            W1024J[600+199] = 16'b0000_0001_0000_0000;
            
            W1024J[700+100] = 16'b0000_0001_0000_0000;
            W1024J[700+101] = 16'b0000_0001_0000_0000;
            W1024J[700+102] = 16'b0000_0001_0000_0000;
            W1024J[700+103] = 16'b0000_0001_0000_0000;
            W1024J[700+104] = 16'b0000_0001_0000_0000;
            W1024J[700+105] = 16'b0000_0001_0000_0000;
            W1024J[700+106] = 16'b0000_0001_0000_0000;
            W1024J[700+107] = 16'b0000_0001_0000_0000;
            W1024J[700+108] = 16'b0000_0001_0000_0000;
            W1024J[700+109] = 16'b0000_0001_0000_0000;
            W1024J[700+110] = 16'b0000_0001_0000_0000;
            W1024J[700+111] = 16'b0000_0001_0000_0000;
            W1024J[700+112] = 16'b0000_0001_0000_0000;
            W1024J[700+113] = 16'b0000_0001_0000_0000;
            W1024J[700+114] = 16'b0000_0001_0000_0000;
            W1024J[700+115] = 16'b0000_0001_0000_0000;
            W1024J[700+116] = 16'b0000_0001_0000_0000;
            W1024J[700+117] = 16'b0000_0001_0000_0000;
            W1024J[700+118] = 16'b0000_0001_0000_0000;
            W1024J[700+119] = 16'b0000_0001_0000_0000;
            W1024J[700+120] = 16'b0000_0001_0000_0000;
            W1024J[700+121] = 16'b0000_0001_0000_0000;
            W1024J[700+122] = 16'b0000_0001_0000_0000;
            W1024J[700+123] = 16'b0000_0001_0000_0000;
            W1024J[700+124] = 16'b0000_0001_0000_0000;
            W1024J[700+125] = 16'b0000_0001_0000_0000;
            W1024J[700+126] = 16'b0000_0001_0000_0000;
            W1024J[700+127] = 16'b0000_0001_0000_0000;
            W1024J[700+128] = 16'b0000_0001_0000_0000;
            W1024J[700+129] = 16'b0000_0001_0000_0000;
            W1024J[700+130] = 16'b0000_0001_0000_0000;
            W1024J[700+131] = 16'b0000_0001_0000_0000;
            W1024J[700+132] = 16'b0000_0001_0000_0000;
            W1024J[700+133] = 16'b0000_0001_0000_0000;
            W1024J[700+134] = 16'b0000_0001_0000_0000;
            W1024J[700+135] = 16'b0000_0001_0000_0000;
            W1024J[700+136] = 16'b0000_0001_0000_0000;
            W1024J[700+137] = 16'b0000_0001_0000_0000;
            W1024J[700+138] = 16'b0000_0001_0000_0000;
            W1024J[700+139] = 16'b0000_0001_0000_0000;
            W1024J[700+140] = 16'b0000_0001_0000_0000;
            W1024J[700+141] = 16'b0000_0001_0000_0000;
            W1024J[700+142] = 16'b0000_0001_0000_0000;
            W1024J[700+143] = 16'b0000_0001_0000_0000;
            W1024J[700+144] = 16'b0000_0001_0000_0000;
            W1024J[700+145] = 16'b0000_0001_0000_0000;
            W1024J[700+146] = 16'b0000_0001_0000_0000;
            W1024J[700+147] = 16'b0000_0001_0000_0000;
            W1024J[700+148] = 16'b0000_0001_0000_0000;
            W1024J[700+149] = 16'b0000_0001_0000_0000;
            W1024J[700+150] = 16'b0000_0001_0000_0000;
            W1024J[700+151] = 16'b0000_0001_0000_0000;
            W1024J[700+152] = 16'b0000_0001_0000_0000;
            W1024J[700+153] = 16'b0000_0001_0000_0000;
            W1024J[700+154] = 16'b0000_0001_0000_0000;
            W1024J[700+155] = 16'b0000_0001_0000_0000;
            W1024J[700+156] = 16'b0000_0001_0000_0000;
            W1024J[700+157] = 16'b0000_0001_0000_0000;
            W1024J[700+158] = 16'b0000_0001_0000_0000;
            W1024J[700+159] = 16'b0000_0001_0000_0000;
            W1024J[700+160] = 16'b0000_0001_0000_0000;
            W1024J[700+161] = 16'b0000_0001_0000_0000;
            W1024J[700+162] = 16'b0000_0001_0000_0000;
            W1024J[700+163] = 16'b0000_0001_0000_0000;
            W1024J[700+164] = 16'b0000_0001_0000_0000;
            W1024J[700+165] = 16'b0000_0001_0000_0000;
            W1024J[700+166] = 16'b0000_0001_0000_0000;
            W1024J[700+167] = 16'b0000_0001_0000_0000;
            W1024J[700+168] = 16'b0000_0001_0000_0000;
            W1024J[700+169] = 16'b0000_0001_0000_0000;
            W1024J[700+170] = 16'b0000_0001_0000_0000;
            W1024J[700+171] = 16'b0000_0001_0000_0000;
            W1024J[700+172] = 16'b0000_0001_0000_0000;
            W1024J[700+173] = 16'b0000_0001_0000_0000;
            W1024J[700+174] = 16'b0000_0001_0000_0000;
            W1024J[700+175] = 16'b0000_0001_0000_0000;
            W1024J[700+176] = 16'b0000_0001_0000_0000;
            W1024J[700+177] = 16'b0000_0001_0000_0000;
            W1024J[700+178] = 16'b0000_0001_0000_0000;
            W1024J[700+179] = 16'b0000_0001_0000_0000;
            W1024J[700+180] = 16'b0000_0001_0000_0000;
            W1024J[700+181] = 16'b0000_0001_0000_0000;
            W1024J[700+182] = 16'b0000_0001_0000_0000;
            W1024J[700+183] = 16'b0000_0001_0000_0000;
            W1024J[700+184] = 16'b0000_0001_0000_0000;
            W1024J[700+185] = 16'b0000_0001_0000_0000;
            W1024J[700+186] = 16'b0000_0001_0000_0000;
            W1024J[700+187] = 16'b0000_0001_0000_0000;
            W1024J[700+188] = 16'b0000_0001_0000_0000;
            W1024J[700+189] = 16'b0000_0001_0000_0000;
            W1024J[700+190] = 16'b0000_0001_0000_0000;
            W1024J[700+191] = 16'b0000_0001_0000_0000;
            W1024J[700+192] = 16'b0000_0001_0000_0000;
            W1024J[700+193] = 16'b0000_0001_0000_0000;
            W1024J[700+194] = 16'b0000_0001_0000_0000;
            W1024J[700+195] = 16'b0000_0001_0000_0000;
            W1024J[700+196] = 16'b0000_0001_0000_0000;
            W1024J[700+197] = 16'b0000_0001_0000_0000;
            W1024J[700+198] = 16'b0000_0001_0000_0000;
            W1024J[700+199] = 16'b0000_0001_0000_0000;
            
            W1024J[800+100] = 16'b0000_0001_0000_0000;
            W1024J[800+101] = 16'b0000_0001_0000_0000;
            W1024J[800+102] = 16'b0000_0001_0000_0000;
            W1024J[800+103] = 16'b0000_0001_0000_0000;
            W1024J[800+104] = 16'b0000_0001_0000_0000;
            W1024J[800+105] = 16'b0000_0001_0000_0000;
            W1024J[800+106] = 16'b0000_0001_0000_0000;
            W1024J[800+107] = 16'b0000_0001_0000_0000;
            W1024J[800+108] = 16'b0000_0001_0000_0000;
            W1024J[800+109] = 16'b0000_0001_0000_0000;
            W1024J[800+110] = 16'b0000_0001_0000_0000;
            W1024J[800+111] = 16'b0000_0001_0000_0000;
            W1024J[800+112] = 16'b0000_0001_0000_0000;
            W1024J[800+113] = 16'b0000_0001_0000_0000;
            W1024J[800+114] = 16'b0000_0001_0000_0000;
            W1024J[800+115] = 16'b0000_0001_0000_0000;
            W1024J[800+116] = 16'b0000_0001_0000_0000;
            W1024J[800+117] = 16'b0000_0001_0000_0000;
            W1024J[800+118] = 16'b0000_0001_0000_0000;
            W1024J[800+119] = 16'b0000_0001_0000_0000;
            W1024J[800+120] = 16'b0000_0001_0000_0000;
            W1024J[800+121] = 16'b0000_0001_0000_0000;
            W1024J[800+122] = 16'b0000_0001_0000_0000;
            W1024J[800+123] = 16'b0000_0001_0000_0000;
            W1024J[800+124] = 16'b0000_0001_0000_0000;
            W1024J[800+125] = 16'b0000_0001_0000_0000;
            W1024J[800+126] = 16'b0000_0001_0000_0000;
            W1024J[800+127] = 16'b0000_0001_0000_0000;
            W1024J[800+128] = 16'b0000_0001_0000_0000;
            W1024J[800+129] = 16'b0000_0001_0000_0000;
            W1024J[800+130] = 16'b0000_0001_0000_0000;
            W1024J[800+131] = 16'b0000_0001_0000_0000;
            W1024J[800+132] = 16'b0000_0001_0000_0000;
            W1024J[800+133] = 16'b0000_0001_0000_0000;
            W1024J[800+134] = 16'b0000_0001_0000_0000;
            W1024J[800+135] = 16'b0000_0001_0000_0000;
            W1024J[800+136] = 16'b0000_0001_0000_0000;
            W1024J[800+137] = 16'b0000_0001_0000_0000;
            W1024J[800+138] = 16'b0000_0001_0000_0000;
            W1024J[800+139] = 16'b0000_0001_0000_0000;
            W1024J[800+140] = 16'b0000_0001_0000_0000;
            W1024J[800+141] = 16'b0000_0001_0000_0000;
            W1024J[800+142] = 16'b0000_0001_0000_0000;
            W1024J[800+143] = 16'b0000_0001_0000_0000;
            W1024J[800+144] = 16'b0000_0001_0000_0000;
            W1024J[800+145] = 16'b0000_0001_0000_0000;
            W1024J[800+146] = 16'b0000_0001_0000_0000;
            W1024J[800+147] = 16'b0000_0001_0000_0000;
            W1024J[800+148] = 16'b0000_0001_0000_0000;
            W1024J[800+149] = 16'b0000_0001_0000_0000;
            W1024J[800+150] = 16'b0000_0001_0000_0000;
            W1024J[800+151] = 16'b0000_0001_0000_0000;
            W1024J[800+152] = 16'b0000_0001_0000_0000;
            W1024J[800+153] = 16'b0000_0001_0000_0000;
            W1024J[800+154] = 16'b0000_0001_0000_0000;
            W1024J[800+155] = 16'b0000_0001_0000_0000;
            W1024J[800+156] = 16'b0000_0001_0000_0000;
            W1024J[800+157] = 16'b0000_0001_0000_0000;
            W1024J[800+158] = 16'b0000_0001_0000_0000;
            W1024J[800+159] = 16'b0000_0001_0000_0000;
            W1024J[800+160] = 16'b0000_0001_0000_0000;
            W1024J[800+161] = 16'b0000_0001_0000_0000;
            W1024J[800+162] = 16'b0000_0001_0000_0000;
            W1024J[800+163] = 16'b0000_0001_0000_0000;
            W1024J[800+164] = 16'b0000_0001_0000_0000;
            W1024J[800+165] = 16'b0000_0001_0000_0000;
            W1024J[800+166] = 16'b0000_0001_0000_0000;
            W1024J[800+167] = 16'b0000_0001_0000_0000;
            W1024J[800+168] = 16'b0000_0001_0000_0000;
            W1024J[800+169] = 16'b0000_0001_0000_0000;
            W1024J[800+170] = 16'b0000_0001_0000_0000;
            W1024J[800+171] = 16'b0000_0001_0000_0000;
            W1024J[800+172] = 16'b0000_0001_0000_0000;
            W1024J[800+173] = 16'b0000_0001_0000_0000;
            W1024J[800+174] = 16'b0000_0001_0000_0000;
            W1024J[800+175] = 16'b0000_0001_0000_0000;
            W1024J[800+176] = 16'b0000_0001_0000_0000;
            W1024J[800+177] = 16'b0000_0001_0000_0000;
            W1024J[800+178] = 16'b0000_0001_0000_0000;
            W1024J[800+179] = 16'b0000_0001_0000_0000;
            W1024J[800+180] = 16'b0000_0001_0000_0000;
            W1024J[800+181] = 16'b0000_0001_0000_0000;
            W1024J[800+182] = 16'b0000_0001_0000_0000;
            W1024J[800+183] = 16'b0000_0001_0000_0000;
            W1024J[800+184] = 16'b0000_0001_0000_0000;
            W1024J[800+185] = 16'b0000_0001_0000_0000;
            W1024J[800+186] = 16'b0000_0001_0000_0000;
            W1024J[800+187] = 16'b0000_0001_0000_0000;
            W1024J[800+188] = 16'b0000_0001_0000_0000;
            W1024J[800+189] = 16'b0000_0001_0000_0000;
            W1024J[800+190] = 16'b0000_0001_0000_0000;
            W1024J[800+191] = 16'b0000_0001_0000_0000;
            W1024J[800+192] = 16'b0000_0001_0000_0000;
            W1024J[800+193] = 16'b0000_0001_0000_0000;
            W1024J[800+194] = 16'b0000_0001_0000_0000;
            W1024J[800+195] = 16'b0000_0001_0000_0000;
            W1024J[800+196] = 16'b0000_0001_0000_0000;
            W1024J[800+197] = 16'b0000_0001_0000_0000;
            W1024J[800+198] = 16'b0000_0001_0000_0000;
            W1024J[800+199] = 16'b0000_0001_0000_0000;
            
            W1024J[1000] = 16'b0000_0001_0000_0000;
            W1024J[1001] = 16'b0000_0001_0000_0000;
            W1024J[1002] = 16'b0000_0001_0000_0000;
            W1024J[1003] = 16'b0000_0001_0000_0000;
            W1024J[1004] = 16'b0000_0001_0000_0000;
            W1024J[1005] = 16'b0000_0001_0000_0000;
            W1024J[1006] = 16'b0000_0001_0000_0000;
            W1024J[1007] = 16'b0000_0001_0000_0000;
            W1024J[1008] = 16'b0000_0001_0000_0000;
            W1024J[1009] = 16'b0000_0001_0000_0000;
            W1024J[1010] = 16'b0000_0001_0000_0000;
            W1024J[1011] = 16'b0000_0001_0000_0000;
            W1024J[1012] = 16'b0000_0001_0000_0000;
            W1024J[1013] = 16'b0000_0001_0000_0000;
            W1024J[1014] = 16'b0000_0001_0000_0000;
            W1024J[1015] = 16'b0000_0001_0000_0000;
            W1024J[1016] = 16'b0000_0001_0000_0000;
            W1024J[1017] = 16'b0000_0001_0000_0000;
            W1024J[1018] = 16'b0000_0001_0000_0000;
            W1024J[1019] = 16'b0000_0001_0000_0000;
            W1024J[1020] = 16'b0000_0001_0000_0000;
            W1024J[1021] = 16'b0000_0001_0000_0000;
            W1024J[1022] = 16'b0000_0001_0000_0000;
            W1024J[1023] = 16'b0000_0001_0000_0000;

            W1024R[0] = 16'b0000000000000000;
W1024R[1] = 16'b1111111111111110;
W1024R[2] = 16'b1111111111111100;
W1024R[3] = 16'b1111111111111011;
W1024R[4] = 16'b1111111111111001;
W1024R[5] = 16'b1111111111111000;
W1024R[6] = 16'b1111111111110110;
W1024R[7] = 16'b1111111111110101;
W1024R[8] = 16'b1111111111110011;
W1024R[9] = 16'b1111111111110001;
W1024R[10] = 16'b1111111111110001;
W1024R[11] = 16'b1111111111110000;
W1024R[12] = 16'b1111111111101110;
W1024R[13] = 16'b1111111111101101;
W1024R[14] = 16'b1111111111101011;
W1024R[15] = 16'b1111111111101010;
W1024R[16] = 16'b1111111111101000;
W1024R[17] = 16'b1111111111100110;
W1024R[18] = 16'b1111111111100101;
W1024R[19] = 16'b1111111111100011;
W1024R[20] = 16'b1111111111100010;
W1024R[21] = 16'b1111111111100000;
W1024R[22] = 16'b1111111111011111;
W1024R[23] = 16'b1111111111011101;
W1024R[24] = 16'b1111111111011011;
W1024R[25] = 16'b1111111111011010;
W1024R[26] = 16'b1111111111011000;
W1024R[27] = 16'b1111111111010111;
W1024R[28] = 16'b1111111111010101;
W1024R[29] = 16'b1111111111010100;
W1024R[30] = 16'b1111111111010010;
W1024R[31] = 16'b1111111111010001;
W1024R[32] = 16'b1111111111001111;
W1024R[33] = 16'b1111111111001110;
W1024R[34] = 16'b1111111111001100;
W1024R[35] = 16'b1111111111001010;
W1024R[36] = 16'b1111111111001001;
W1024R[37] = 16'b1111111111000111;
W1024R[38] = 16'b1111111111000110;
W1024R[39] = 16'b1111111111000100;
W1024R[40] = 16'b1111111111000011;
W1024R[41] = 16'b1111111111000001;
W1024R[42] = 16'b1111111111000000;
W1024R[43] = 16'b1111111110111110;
W1024R[44] = 16'b1111111110111101;
W1024R[45] = 16'b1111111110111011;
W1024R[46] = 16'b1111111110111010;
W1024R[47] = 16'b1111111110111000;
W1024R[48] = 16'b1111111110110111;
W1024R[49] = 16'b1111111110110101;
W1024R[50] = 16'b1111111110110100;
W1024R[51] = 16'b1111111110110010;
W1024R[52] = 16'b1111111110110001;
W1024R[53] = 16'b1111111110101111;
W1024R[54] = 16'b1111111110101110;
W1024R[55] = 16'b1111111110101100;
W1024R[56] = 16'b1111111110101011;
W1024R[57] = 16'b1111111110101001;
W1024R[58] = 16'b1111111110101000;
W1024R[59] = 16'b1111111110100110;
W1024R[60] = 16'b1111111110100101;
W1024R[61] = 16'b1111111110100011;
W1024R[62] = 16'b1111111110100010;
W1024R[63] = 16'b1111111110100000;
W1024R[64] = 16'b1111111110011111;
W1024R[65] = 16'b1111111110011110;
W1024R[66] = 16'b1111111110011100;
W1024R[67] = 16'b1111111110011011;
W1024R[68] = 16'b1111111110011001;
W1024R[69] = 16'b1111111110011000;
W1024R[70] = 16'b1111111110010110;
W1024R[71] = 16'b1111111110010101;
W1024R[72] = 16'b1111111110010011;
W1024R[73] = 16'b1111111110010010;
W1024R[74] = 16'b1111111110010001;
W1024R[75] = 16'b1111111110001111;
W1024R[76] = 16'b1111111110001110;
W1024R[77] = 16'b1111111110001100;
W1024R[78] = 16'b1111111110001011;
W1024R[79] = 16'b1111111110001010;
W1024R[80] = 16'b1111111110001000;
W1024R[81] = 16'b1111111110000111;
W1024R[82] = 16'b1111111110000101;
W1024R[83] = 16'b1111111110000100;
W1024R[84] = 16'b1111111110000011;
W1024R[85] = 16'b1111111110000001;
W1024R[86] = 16'b1111111110000000;
W1024R[87] = 16'b1111111101111111;
W1024R[88] = 16'b1111111101111101;
W1024R[89] = 16'b1111111101111100;
W1024R[90] = 16'b1111111101111011;
W1024R[91] = 16'b1111111101111001;
W1024R[92] = 16'b1111111101111000;
W1024R[93] = 16'b1111111101110111;
W1024R[94] = 16'b1111111101110101;
W1024R[95] = 16'b1111111101110100;
W1024R[96] = 16'b1111111101110011;
W1024R[97] = 16'b1111111101110001;
W1024R[98] = 16'b1111111101110000;
W1024R[99] = 16'b1111111101101111;

W1024R[100] = 16'b1111111101101100;
W1024R[101] = 16'b1111111101101100;
W1024R[102] = 16'b1111111101101011;
W1024R[103] = 16'b1111111101101010;
W1024R[104] = 16'b1111111101101000;
W1024R[105] = 16'b1111111101100111;
W1024R[106] = 16'b1111111101100110;
W1024R[107] = 16'b1111111101100100;
W1024R[108] = 16'b1111111101100011;
W1024R[109] = 16'b1111111101100010;
W1024R[110] = 16'b1111111101100001;
W1024R[111] = 16'b1111111101100000;
W1024R[112] = 16'b1111111101011101;
W1024R[113] = 16'b1111111101011100;
W1024R[114] = 16'b1111111101011011;
W1024R[115] = 16'b1111111101011001;
W1024R[116] = 16'b1111111101011000;
W1024R[117] = 16'b1111111101010111;
W1024R[118] = 16'b1111111101010110;
W1024R[119] = 16'b1111111101010101;
W1024R[120] = 16'b1111111101010100;
W1024R[121] = 16'b1111111101010010;
W1024R[122] = 16'b1111111101010001;
W1024R[123] = 16'b1111111101010000;
W1024R[124] = 16'b1111111101001111;
W1024R[125] = 16'b1111111101001110;
W1024R[126] = 16'b1111111101001101;
W1024R[127] = 16'b1111111101001100;
W1024R[128] = 16'b1111111101001010;
W1024R[129] = 16'b1111111101001001;
W1024R[130] = 16'b1111111101001000;
W1024R[131] = 16'b1111111101000111;
W1024R[132] = 16'b1111111101000110;
W1024R[133] = 16'b1111111101000101;
W1024R[134] = 16'b1111111101000100;
W1024R[135] = 16'b1111111101000011;
W1024R[136] = 16'b1111111101000010;
W1024R[137] = 16'b1111111101000001;
W1024R[138] = 16'b1111111101000000;
W1024R[139] = 16'b1111111100111111;
W1024R[140] = 16'b1111111100111110;
W1024R[141] = 16'b1111111100111101;
W1024R[142] = 16'b1111111100111100;
W1024R[143] = 16'b1111111100111011;
W1024R[144] = 16'b1111111100111010;
W1024R[145] = 16'b1111111100111001;
W1024R[146] = 16'b1111111100111000;
W1024R[147] = 16'b1111111100110111;
W1024R[148] = 16'b1111111100110110;
W1024R[149] = 16'b1111111100110101;
W1024R[150] = 16'b1111111100110100;
W1024R[151] = 16'b1111111100110011;
W1024R[152] = 16'b1111111100110010;
W1024R[153] = 16'b1111111100110001;
W1024R[154] = 16'b1111111100110000;
W1024R[155] = 16'b1111111100101111;
W1024R[156] = 16'b1111111100101110;
W1024R[157] = 16'b1111111100101101;
W1024R[158] = 16'b1111111100101100;
W1024R[159] = 16'b1111111100101100;
W1024R[160] = 16'b1111111100101011;
W1024R[161] = 16'b1111111100101010;
W1024R[162] = 16'b1111111100101001;
W1024R[163] = 16'b1111111100101000;
W1024R[164] = 16'b1111111100100111;
W1024R[165] = 16'b1111111100100110;
W1024R[166] = 16'b1111111100100110;
W1024R[167] = 16'b1111111100100101;
W1024R[168] = 16'b1111111100100100;
W1024R[169] = 16'b1111111100100011;
W1024R[170] = 16'b1111111100100010;
W1024R[171] = 16'b1111111100100010;
W1024R[172] = 16'b1111111100100001;
W1024R[173] = 16'b1111111100100000;
W1024R[174] = 16'b1111111100011111;
W1024R[175] = 16'b1111111100011110;
W1024R[176] = 16'b1111111100011110;
W1024R[177] = 16'b1111111100011101;
W1024R[178] = 16'b1111111100011100;
W1024R[179] = 16'b1111111100011100;
W1024R[180] = 16'b1111111100011011;
W1024R[181] = 16'b1111111100011010;
W1024R[182] = 16'b1111111100011001;
W1024R[183] = 16'b1111111100011001;
W1024R[184] = 16'b1111111100011000;
W1024R[185] = 16'b1111111100010111;
W1024R[186] = 16'b1111111100010111;
W1024R[187] = 16'b1111111100010110;
W1024R[188] = 16'b1111111100010101;
W1024R[189] = 16'b1111111100010101;
W1024R[190] = 16'b1111111100010100;
W1024R[191] = 16'b1111111100010100;
W1024R[192] = 16'b1111111100010011;
W1024R[193] = 16'b1111111100010010;
W1024R[194] = 16'b1111111100010010;
W1024R[195] = 16'b1111111100010010;
W1024R[196] = 16'b1111111100010001;
W1024R[197] = 16'b1111111100010001;
W1024R[198] = 16'b1111111100010000;
W1024R[199] = 16'b1111111100010000;

W1024R[100+100] = 16'b1111111100001110;
W1024R[100+101] = 16'b1111111100001110;
W1024R[100+102] = 16'b1111111100001101;
W1024R[100+103] = 16'b1111111100001101;
W1024R[100+104] = 16'b1111111100001100;
W1024R[100+105] = 16'b1111111100001100;
W1024R[100+106] = 16'b1111111100001011;
W1024R[100+107] = 16'b1111111100001011;
W1024R[100+108] = 16'b1111111100001011;
W1024R[100+109] = 16'b1111111100001010;
W1024R[100+110] = 16'b1111111100001010;
W1024R[100+111] = 16'b1111111100001001;
W1024R[100+112] = 16'b1111111100001001;
W1024R[100+113] = 16'b1111111100001000;
W1024R[100+114] = 16'b1111111100001000;
W1024R[100+115] = 16'b1111111100001000;
W1024R[100+116] = 16'b1111111100000111;
W1024R[100+117] = 16'b1111111100000111;
W1024R[100+118] = 16'b1111111100000110;
W1024R[100+119] = 16'b1111111100000110;
W1024R[100+120] = 16'b1111111100000110;
W1024R[100+121] = 16'b1111111100000101;
W1024R[100+122] = 16'b1111111100000101;
W1024R[100+123] = 16'b1111111100000101;
W1024R[100+124] = 16'b1111111100000100;
W1024R[100+125] = 16'b1111111100000100;
W1024R[100+126] = 16'b1111111100000100;
W1024R[100+127] = 16'b1111111100000100;
W1024R[100+128] = 16'b1111111100000011;
W1024R[100+129] = 16'b1111111100000011;
W1024R[100+130] = 16'b1111111100000011;
W1024R[100+131] = 16'b1111111100000011;
W1024R[100+132] = 16'b1111111100000010;
W1024R[100+133] = 16'b1111111100000010;
W1024R[100+134] = 16'b1111111100000010;
W1024R[100+135] = 16'b1111111100000010;
W1024R[100+136] = 16'b1111111100000001;
W1024R[100+137] = 16'b1111111100000001;
W1024R[100+138] = 16'b1111111100000001;
W1024R[100+139] = 16'b1111111100000001;
W1024R[100+140] = 16'b1111111100000001;
W1024R[100+141] = 16'b1111111100000001;
W1024R[100+142] = 16'b1111111100000001;
W1024R[100+143] = 16'b1111111100000000;
W1024R[100+144] = 16'b1111111100000000;
W1024R[100+145] = 16'b1111111100000000;
W1024R[100+146] = 16'b1111111100000000;
W1024R[100+147] = 16'b1111111100000000;
W1024R[100+148] = 16'b1111111100000000;
W1024R[100+149] = 16'b1111111100000000;
W1024R[100+150] = 16'b1111111100000000;
W1024R[100+151] = 16'b1111111100000000;
W1024R[100+152] = 16'b1111111100000000;
W1024R[100+153] = 16'b1111111100000000;
W1024R[100+154] = 16'b1111111100000000;
W1024R[100+155] = 16'b1111111100000000;
W1024R[100+156] = 16'b1111111100000000;
W1024R[100+157] = 16'b1111111100000000;
W1024R[100+158] = 16'b1111111100000000;
W1024R[100+159] = 16'b1111111100000000;
W1024R[100+160] = 16'b1111111100000000;
W1024R[100+161] = 16'b1111111100000000;
W1024R[100+162] = 16'b1111111100000000;
W1024R[100+163] = 16'b1111111100000000;
W1024R[100+164] = 16'b1111111100000000;
W1024R[100+165] = 16'b1111111100000000;
W1024R[100+166] = 16'b1111111100000000;
W1024R[100+167] = 16'b1111111100000000;
W1024R[100+168] = 16'b1111111100000000;
W1024R[100+169] = 16'b1111111100000000;
W1024R[100+170] = 16'b1111111100000000;
W1024R[100+171] = 16'b1111111100000000;
W1024R[100+172] = 16'b1111111100000001;
W1024R[100+173] = 16'b1111111100000001;
W1024R[100+174] = 16'b1111111100000001;
W1024R[100+175] = 16'b1111111100000001;
W1024R[100+176] = 16'b1111111100000001;
W1024R[100+177] = 16'b1111111100000001;
W1024R[100+178] = 16'b1111111100000010;
W1024R[100+179] = 16'b1111111100000010;
W1024R[100+180] = 16'b1111111100000010;
W1024R[100+181] = 16'b1111111100000010;
W1024R[100+182] = 16'b1111111100000011;
W1024R[100+183] = 16'b1111111100000011;
W1024R[100+184] = 16'b1111111100000011;
W1024R[100+185] = 16'b1111111100000011;
W1024R[100+186] = 16'b1111111100000100;
W1024R[100+187] = 16'b1111111100000100;
W1024R[100+188] = 16'b1111111100000100;
W1024R[100+189] = 16'b1111111100000100;
W1024R[100+190] = 16'b1111111100000101;
W1024R[100+191] = 16'b1111111100000101;
W1024R[100+192] = 16'b1111111100000101;
W1024R[100+193] = 16'b1111111100000110;
W1024R[100+194] = 16'b1111111100000110;
W1024R[100+195] = 16'b1111111100000110;
W1024R[100+196] = 16'b1111111100000111;
W1024R[100+197] = 16'b1111111100000111;
W1024R[100+198] = 16'b1111111100001000;
W1024R[100+199] = 16'b1111111100001000;



W1024R[200+100] = 16'b1111111100001001;
W1024R[200+101] = 16'b1111111100001001;
W1024R[200+102] = 16'b1111111100001010;
W1024R[200+103] = 16'b1111111100001010;
W1024R[200+104] = 16'b1111111100001011;
W1024R[200+105] = 16'b1111111100001011;
W1024R[200+106] = 16'b1111111100001011;
W1024R[200+107] = 16'b1111111100001100;
W1024R[200+108] = 16'b1111111100001100;
W1024R[200+109] = 16'b1111111100001101;
W1024R[200+110] = 16'b1111111100001101;
W1024R[200+111] = 16'b1111111100001110;
W1024R[200+112] = 16'b1111111100001110;
W1024R[200+113] = 16'b1111111100001111;
W1024R[200+114] = 16'b1111111100010000;
W1024R[200+115] = 16'b1111111100010000;
W1024R[200+116] = 16'b1111111100010001;
W1024R[200+117] = 16'b1111111100010001;
W1024R[200+118] = 16'b1111111100010010;
W1024R[200+119] = 16'b1111111100010010;
W1024R[200+120] = 16'b1111111100010011;
W1024R[200+121] = 16'b1111111100010100;
W1024R[200+122] = 16'b1111111100010100;
W1024R[200+123] = 16'b1111111100010101;
W1024R[200+124] = 16'b1111111100010101;
W1024R[200+125] = 16'b1111111100010110;
W1024R[200+126] = 16'b1111111100010111;
W1024R[200+127] = 16'b1111111100010111;
W1024R[200+128] = 16'b1111111100011000;
W1024R[200+129] = 16'b1111111100011001;
W1024R[200+130] = 16'b1111111100011001;
W1024R[200+131] = 16'b1111111100011010;
W1024R[200+132] = 16'b1111111100011011;
W1024R[200+133] = 16'b1111111100011100;
W1024R[200+134] = 16'b1111111100011100;
W1024R[200+135] = 16'b1111111100011101;
W1024R[200+136] = 16'b1111111100011110;
W1024R[200+137] = 16'b1111111100011110;
W1024R[200+138] = 16'b1111111100011111;
W1024R[200+139] = 16'b1111111100100000;
W1024R[200+140] = 16'b1111111100100001;
W1024R[200+141] = 16'b1111111100100010;
W1024R[200+142] = 16'b1111111100100010;
W1024R[200+143] = 16'b1111111100100011;
W1024R[200+144] = 16'b1111111100100100;
W1024R[200+145] = 16'b1111111100100101;
W1024R[200+146] = 16'b1111111100100110;
W1024R[200+147] = 16'b1111111100100110;
W1024R[200+148] = 16'b1111111100100111;
W1024R[200+149] = 16'b1111111100100110;
W1024R[200+150] = 16'b1111111100100111;
W1024R[200+151] = 16'b1111111100101000;
W1024R[200+152] = 16'b1111111100101001;
W1024R[200+153] = 16'b1111111100101010;
W1024R[200+154] = 16'b1111111100101011;
W1024R[200+155] = 16'b1111111100101100;
W1024R[200+156] = 16'b1111111100101100;
W1024R[200+157] = 16'b1111111100101101;
W1024R[200+158] = 16'b1111111100101110;
W1024R[200+159] = 16'b1111111100101111;
W1024R[200+160] = 16'b1111111100110000;
W1024R[200+161] = 16'b1111111100110001;
W1024R[200+162] = 16'b1111111100110010;
W1024R[200+163] = 16'b1111111100110011;
W1024R[200+164] = 16'b1111111100110100;
W1024R[200+165] = 16'b1111111100110101;
W1024R[200+166] = 16'b1111111100110111;
W1024R[200+167] = 16'b1111111100111000;
W1024R[200+168] = 16'b1111111100111001;
W1024R[200+169] = 16'b1111111100111010;
W1024R[200+170] = 16'b1111111100111011;
W1024R[200+171] = 16'b1111111100111100;
W1024R[200+172] = 16'b1111111100111101;
W1024R[200+173] = 16'b1111111100111110;
W1024R[200+174] = 16'b1111111100111111;
W1024R[200+175] = 16'b1111111101000000;
W1024R[200+176] = 16'b1111111101000001;
W1024R[200+177] = 16'b1111111101000010;
W1024R[200+178] = 16'b1111111101000011;
W1024R[200+179] = 16'b1111111101000100;
W1024R[200+180] = 16'b1111111101000101;
W1024R[200+181] = 16'b1111111101000110;
W1024R[200+182] = 16'b1111111101000111;
W1024R[200+183] = 16'b1111111101001000;
W1024R[200+184] = 16'b1111111101001001;
W1024R[200+185] = 16'b1111111101001010;
W1024R[200+186] = 16'b1111111101001100;
W1024R[200+187] = 16'b1111111101001101;
W1024R[200+188] = 16'b1111111101001110;
W1024R[200+189] = 16'b1111111101001111;
W1024R[200+190] = 16'b1111111101010000;
W1024R[200+191] = 16'b1111111101010001;
W1024R[200+192] = 16'b1111111101010010;
W1024R[200+193] = 16'b1111111101010100;
W1024R[200+194] = 16'b1111111101010101;
W1024R[200+195] = 16'b1111111101010110;
W1024R[200+196] = 16'b1111111101010111;
W1024R[200+197] = 16'b1111111101011000;
W1024R[200+198] = 16'b1111111101011001;
W1024R[200+199] = 16'b1111111101011011;

W1024R[300+100] = 16'b0000_0001_0000_0000;
W1024R[300+101] = 16'b0000_0001_0000_0000;
W1024R[300+102] = 16'b0000_0001_0000_0000;
W1024R[300+103] = 16'b0000_0001_0000_0000;
W1024R[300+104] = 16'b0000_0001_0000_0000;
W1024R[300+105] = 16'b0000_0001_0000_0000;
W1024R[300+106] = 16'b0000_0001_0000_0000;
W1024R[300+107] = 16'b0000_0001_0000_0000;
W1024R[300+108] = 16'b0000_0001_0000_0000;
W1024R[300+109] = 16'b0000_0001_0000_0000;
W1024R[300+110] = 16'b0000_0001_0000_0000;
W1024R[300+111] = 16'b0000_0001_0000_0000;
W1024R[300+112] = 16'b0000_0001_0000_0000;
W1024R[300+113] = 16'b0000_0001_0000_0000;
W1024R[300+114] = 16'b0000_0001_0000_0000;
W1024R[300+115] = 16'b0000_0001_0000_0000;
W1024R[300+116] = 16'b0000_0001_0000_0000;
W1024R[300+117] = 16'b0000_0001_0000_0000;
W1024R[300+118] = 16'b0000_0001_0000_0000;
W1024R[300+119] = 16'b0000_0001_0000_0000;
W1024R[300+120] = 16'b0000_0001_0000_0000;
W1024R[300+121] = 16'b0000_0001_0000_0000;
W1024R[300+122] = 16'b0000_0001_0000_0000;
W1024R[300+123] = 16'b0000_0001_0000_0000;
W1024R[300+124] = 16'b0000_0001_0000_0000;
W1024R[300+125] = 16'b0000_0001_0000_0000;
W1024R[300+126] = 16'b0000_0001_0000_0000;
W1024R[300+127] = 16'b0000_0001_0000_0000;
W1024R[300+128] = 16'b0000_0001_0000_0000;
W1024R[300+129] = 16'b0000_0001_0000_0000;
W1024R[300+130] = 16'b0000_0001_0000_0000;
W1024R[300+131] = 16'b0000_0001_0000_0000;
W1024R[300+132] = 16'b0000_0001_0000_0000;
W1024R[300+133] = 16'b0000_0001_0000_0000;
W1024R[300+134] = 16'b0000_0001_0000_0000;
W1024R[300+135] = 16'b0000_0001_0000_0000;
W1024R[300+136] = 16'b0000_0001_0000_0000;
W1024R[300+137] = 16'b0000_0001_0000_0000;
W1024R[300+138] = 16'b0000_0001_0000_0000;
W1024R[300+139] = 16'b0000_0001_0000_0000;
W1024R[300+140] = 16'b0000_0001_0000_0000;
W1024R[300+141] = 16'b0000_0001_0000_0000;
W1024R[300+142] = 16'b0000_0001_0000_0000;
W1024R[300+143] = 16'b0000_0001_0000_0000;
W1024R[300+144] = 16'b0000_0001_0000_0000;
W1024R[300+145] = 16'b0000_0001_0000_0000;
W1024R[300+146] = 16'b0000_0001_0000_0000;
W1024R[300+147] = 16'b0000_0001_0000_0000;
W1024R[300+148] = 16'b0000_0001_0000_0000;
W1024R[300+149] = 16'b0000_0001_0000_0000;
W1024R[300+150] = 16'b0000_0001_0000_0000;
W1024R[300+151] = 16'b0000_0001_0000_0000;
W1024R[300+152] = 16'b0000_0001_0000_0000;
W1024R[300+153] = 16'b0000_0001_0000_0000;
W1024R[300+154] = 16'b0000_0001_0000_0000;
W1024R[300+155] = 16'b0000_0001_0000_0000;
W1024R[300+156] = 16'b0000_0001_0000_0000;
W1024R[300+157] = 16'b0000_0001_0000_0000;
W1024R[300+158] = 16'b0000_0001_0000_0000;
W1024R[300+159] = 16'b0000_0001_0000_0000;
W1024R[300+160] = 16'b0000_0001_0000_0000;
W1024R[300+161] = 16'b0000_0001_0000_0000;
W1024R[300+162] = 16'b0000_0001_0000_0000;
W1024R[300+163] = 16'b0000_0001_0000_0000;
W1024R[300+164] = 16'b0000_0001_0000_0000;
W1024R[300+165] = 16'b0000_0001_0000_0000;
W1024R[300+166] = 16'b0000_0001_0000_0000;
W1024R[300+167] = 16'b0000_0001_0000_0000;
W1024R[300+168] = 16'b0000_0001_0000_0000;
W1024R[300+169] = 16'b0000_0001_0000_0000;
W1024R[300+170] = 16'b0000_0001_0000_0000;
W1024R[300+171] = 16'b0000_0001_0000_0000;
W1024R[300+172] = 16'b0000_0001_0000_0000;
W1024R[300+173] = 16'b0000_0001_0000_0000;
W1024R[300+174] = 16'b0000_0001_0000_0000;
W1024R[300+175] = 16'b0000_0001_0000_0000;
W1024R[300+176] = 16'b0000_0001_0000_0000;
W1024R[300+177] = 16'b0000_0001_0000_0000;
W1024R[300+178] = 16'b0000_0001_0000_0000;
W1024R[300+179] = 16'b0000_0001_0000_0000;
W1024R[300+180] = 16'b0000_0001_0000_0000;
W1024R[300+181] = 16'b0000_0001_0000_0000;
W1024R[300+182] = 16'b0000_0001_0000_0000;
W1024R[300+183] = 16'b0000_0001_0000_0000;
W1024R[300+184] = 16'b0000_0001_0000_0000;
W1024R[300+185] = 16'b0000_0001_0000_0000;
W1024R[300+186] = 16'b0000_0001_0000_0000;
W1024R[300+187] = 16'b0000_0001_0000_0000;
W1024R[300+188] = 16'b0000_0001_0000_0000;
W1024R[300+189] = 16'b0000_0001_0000_0000;
W1024R[300+190] = 16'b0000_0001_0000_0000;
W1024R[300+191] = 16'b0000_0001_0000_0000;
W1024R[300+192] = 16'b0000_0001_0000_0000;
W1024R[300+193] = 16'b0000_0001_0000_0000;
W1024R[300+194] = 16'b0000_0001_0000_0000;
W1024R[300+195] = 16'b0000_0001_0000_0000;
W1024R[300+196] = 16'b0000_0001_0000_0000;
W1024R[300+197] = 16'b0000_0001_0000_0000;
W1024R[300+198] = 16'b0000_0001_0000_0000;
W1024R[300+199] = 16'b0000_0001_0000_0000;

W1024R[400+100] = 16'b0000_0001_0000_0000;
W1024R[400+101] = 16'b0000_0001_0000_0000;
W1024R[400+102] = 16'b0000_0001_0000_0000;
W1024R[400+103] = 16'b0000_0001_0000_0000;
W1024R[400+104] = 16'b0000_0001_0000_0000;
W1024R[400+105] = 16'b0000_0001_0000_0000;
W1024R[400+106] = 16'b0000_0001_0000_0000;
W1024R[400+107] = 16'b0000_0001_0000_0000;
W1024R[400+108] = 16'b0000_0001_0000_0000;
W1024R[400+109] = 16'b0000_0001_0000_0000;
W1024R[400+110] = 16'b0000_0001_0000_0000;
W1024R[400+111] = 16'b0000_0001_0000_0000;
W1024R[400+112] = 16'b0000_0001_0000_0000;



W1024R[400+113] = 16'b0000_0001_0000_0000;
W1024R[400+114] = 16'b0000_0001_0000_0000;
W1024R[400+115] = 16'b0000_0001_0000_0000;
W1024R[400+116] = 16'b0000_0001_0000_0000;
W1024R[400+117] = 16'b0000_0001_0000_0000;
W1024R[400+118] = 16'b0000_0001_0000_0000;
W1024R[400+119] = 16'b0000_0001_0000_0000;
W1024R[400+120] = 16'b0000_0001_0000_0000;
W1024R[400+121] = 16'b0000_0001_0000_0000;
W1024R[400+122] = 16'b0000_0001_0000_0000;
W1024R[400+123] = 16'b0000_0001_0000_0000;
W1024R[400+124] = 16'b0000_0001_0000_0000;
W1024R[400+125] = 16'b0000_0001_0000_0000;
W1024R[400+126] = 16'b0000_0001_0000_0000;
W1024R[400+127] = 16'b0000_0001_0000_0000;
W1024R[400+128] = 16'b0000_0001_0000_0000;
W1024R[400+129] = 16'b0000_0001_0000_0000;
W1024R[400+130] = 16'b0000_0001_0000_0000;
W1024R[400+131] = 16'b0000_0001_0000_0000;
W1024R[400+132] = 16'b0000_0001_0000_0000;
W1024R[400+133] = 16'b0000_0001_0000_0000;
W1024R[400+134] = 16'b0000_0001_0000_0000;
W1024R[400+135] = 16'b0000_0001_0000_0000;
W1024R[400+136] = 16'b0000_0001_0000_0000;
W1024R[400+137] = 16'b0000_0001_0000_0000;
W1024R[400+138] = 16'b0000_0001_0000_0000;
W1024R[400+139] = 16'b0000_0001_0000_0000;
W1024R[400+140] = 16'b0000_0001_0000_0000;
W1024R[400+141] = 16'b0000_0001_0000_0000;
W1024R[400+142] = 16'b0000_0001_0000_0000;
W1024R[400+143] = 16'b0000_0001_0000_0000;
W1024R[400+144] = 16'b0000_0001_0000_0000;
W1024R[400+145] = 16'b0000_0001_0000_0000;
W1024R[400+146] = 16'b0000_0001_0000_0000;
W1024R[400+147] = 16'b0000_0001_0000_0000;
W1024R[400+148] = 16'b0000_0001_0000_0000;
W1024R[400+149] = 16'b0000_0001_0000_0000;
W1024R[400+150] = 16'b0000_0001_0000_0000;
W1024R[400+151] = 16'b0000_0001_0000_0000;
W1024R[400+152] = 16'b0000_0001_0000_0000;
W1024R[400+153] = 16'b0000_0001_0000_0000;
W1024R[400+154] = 16'b0000_0001_0000_0000;
W1024R[400+155] = 16'b0000_0001_0000_0000;
W1024R[400+156] = 16'b0000_0001_0000_0000;
W1024R[400+157] = 16'b0000_0001_0000_0000;
W1024R[400+158] = 16'b0000_0001_0000_0000;
W1024R[400+159] = 16'b0000_0001_0000_0000;
W1024R[400+160] = 16'b0000_0001_0000_0000;
W1024R[400+161] = 16'b0000_0001_0000_0000;
W1024R[400+162] = 16'b0000_0001_0000_0000;
W1024R[400+163] = 16'b0000_0001_0000_0000;
W1024R[400+164] = 16'b0000_0001_0000_0000;
W1024R[400+165] = 16'b0000_0001_0000_0000;
W1024R[400+166] = 16'b0000_0001_0000_0000;
W1024R[400+167] = 16'b0000_0001_0000_0000;
W1024R[400+168] = 16'b0000_0001_0000_0000;
W1024R[400+169] = 16'b0000_0001_0000_0000;
W1024R[400+170] = 16'b0000_0001_0000_0000;
W1024R[400+171] = 16'b0000_0001_0000_0000;
W1024R[400+172] = 16'b0000_0001_0000_0000;
W1024R[400+173] = 16'b0000_0001_0000_0000;
W1024R[400+174] = 16'b0000_0001_0000_0000;
W1024R[400+175] = 16'b0000_0001_0000_0000;
W1024R[400+176] = 16'b0000_0001_0000_0000;
W1024R[400+177] = 16'b0000_0001_0000_0000;
W1024R[400+178] = 16'b0000_0001_0000_0000;
W1024R[400+179] = 16'b0000_0001_0000_0000;
W1024R[400+180] = 16'b0000_0001_0000_0000;
W1024R[400+181] = 16'b0000_0001_0000_0000;
W1024R[400+182] = 16'b0000_0001_0000_0000;
W1024R[400+183] = 16'b0000_0001_0000_0000;
W1024R[400+184] = 16'b0000_0001_0000_0000;
W1024R[400+185] = 16'b0000_0001_0000_0000;
W1024R[400+186] = 16'b0000_0001_0000_0000;
W1024R[400+187] = 16'b0000_0001_0000_0000;
W1024R[400+188] = 16'b0000_0001_0000_0000;
W1024R[400+189] = 16'b0000_0001_0000_0000;
W1024R[400+190] = 16'b0000_0001_0000_0000;
W1024R[400+191] = 16'b0000_0001_0000_0000;
W1024R[400+192] = 16'b0000_0001_0000_0000;
W1024R[400+193] = 16'b0000_0001_0000_0000;
W1024R[400+194] = 16'b0000_0001_0000_0000;
W1024R[400+195] = 16'b0000_0001_0000_0000;
W1024R[400+196] = 16'b0000_0001_0000_0000;
W1024R[400+197] = 16'b0000_0001_0000_0000;
W1024R[400+198] = 16'b0000_0001_0000_0000;
W1024R[400+199] = 16'b0000_0001_0000_0000;

W1024R[500+100] = 16'b0000_0001_0000_0000;
W1024R[500+101] = 16'b0000_0001_0000_0000;
W1024R[500+102] = 16'b0000_0001_0000_0000;
W1024R[500+103] = 16'b0000_0001_0000_0000;
W1024R[500+104] = 16'b0000_0001_0000_0000;
W1024R[500+105] = 16'b0000_0001_0000_0000;
W1024R[500+106] = 16'b0000_0001_0000_0000;
W1024R[500+107] = 16'b0000_0001_0000_0000;
W1024R[500+108] = 16'b0000_0001_0000_0000;
W1024R[500+109] = 16'b0000_0001_0000_0000;
W1024R[500+110] = 16'b0000_0001_0000_0000;
W1024R[500+111] = 16'b0000_0001_0000_0000;
W1024R[500+112] = 16'b0000_0001_0000_0000;
W1024R[500+113] = 16'b0000_0001_0000_0000;
W1024R[500+114] = 16'b0000_0001_0000_0000;
W1024R[500+115] = 16'b0000_0001_0000_0000;
W1024R[500+116] = 16'b0000_0001_0000_0000;
W1024R[500+117] = 16'b0000_0001_0000_0000;
W1024R[500+118] = 16'b0000_0001_0000_0000;
W1024R[500+119] = 16'b0000_0001_0000_0000;
W1024R[500+120] = 16'b0000_0001_0000_0000;
W1024R[500+121] = 16'b0000_0001_0000_0000;
W1024R[500+122] = 16'b0000_0001_0000_0000;
W1024R[500+123] = 16'b0000_0001_0000_0000;
W1024R[500+124] = 16'b0000_0001_0000_0000;
W1024R[500+125] = 16'b0000_0001_0000_0000;
W1024R[500+126] = 16'b0000_0001_0000_0000;
W1024R[500+127] = 16'b0000_0001_0000_0000;
W1024R[500+128] = 16'b0000_0001_0000_0000;
W1024R[500+129] = 16'b0000_0001_0000_0000;
W1024R[500+130] = 16'b0000_0001_0000_0000;
W1024R[500+131] = 16'b0000_0001_0000_0000;
W1024R[500+132] = 16'b0000_0001_0000_0000;
W1024R[500+133] = 16'b0000_0001_0000_0000;
W1024R[500+134] = 16'b0000_0001_0000_0000;
W1024R[500+135] = 16'b0000_0001_0000_0000;
W1024R[500+136] = 16'b0000_0001_0000_0000;
W1024R[500+137] = 16'b0000_0001_0000_0000;
W1024R[500+138] = 16'b0000_0001_0000_0000;
W1024R[500+139] = 16'b0000_0001_0000_0000;
W1024R[500+140] = 16'b0000_0001_0000_0000;
W1024R[500+141] = 16'b0000_0001_0000_0000;
W1024R[500+142] = 16'b0000_0001_0000_0000;
W1024R[500+143] = 16'b0000_0001_0000_0000;
W1024R[500+144] = 16'b0000_0001_0000_0000;
W1024R[500+145] = 16'b0000_0001_0000_0000;
W1024R[500+146] = 16'b0000_0001_0000_0000;
W1024R[500+147] = 16'b0000_0001_0000_0000;
W1024R[500+148] = 16'b0000_0001_0000_0000;
W1024R[500+149] = 16'b0000_0001_0000_0000;
W1024R[500+150] = 16'b0000_0001_0000_0000;
W1024R[500+151] = 16'b0000_0001_0000_0000;
W1024R[500+152] = 16'b0000_0001_0000_0000;
W1024R[500+153] = 16'b0000_0001_0000_0000;
W1024R[500+154] = 16'b0000_0001_0000_0000;
W1024R[500+155] = 16'b0000_0001_0000_0000;
W1024R[500+156] = 16'b0000_0001_0000_0000;
W1024R[500+157] = 16'b0000_0001_0000_0000;
W1024R[500+158] = 16'b0000_0001_0000_0000;
W1024R[500+159] = 16'b0000_0001_0000_0000;
W1024R[500+160] = 16'b0000_0001_0000_0000;
W1024R[500+161] = 16'b0000_0001_0000_0000;
W1024R[500+162] = 16'b0000_0001_0000_0000;
W1024R[500+163] = 16'b0000_0001_0000_0000;
W1024R[500+164] = 16'b0000_0001_0000_0000;
W1024R[500+165] = 16'b0000_0001_0000_0000;
W1024R[500+166] = 16'b0000_0001_0000_0000;
W1024R[500+167] = 16'b0000_0001_0000_0000;
W1024R[500+168] = 16'b0000_0001_0000_0000;
W1024R[500+169] = 16'b0000_0001_0000_0000;
W1024R[500+170] = 16'b0000_0001_0000_0000;
W1024R[500+171] = 16'b0000_0001_0000_0000;
W1024R[500+172] = 16'b0000_0001_0000_0000;
W1024R[500+173] = 16'b0000_0001_0000_0000;
W1024R[500+174] = 16'b0000_0001_0000_0000;
W1024R[500+175] = 16'b0000_0001_0000_0000;
W1024R[500+176] = 16'b0000_0001_0000_0000;
W1024R[500+177] = 16'b0000_0001_0000_0000;
W1024R[500+178] = 16'b0000_0001_0000_0000;
W1024R[500+179] = 16'b0000_0001_0000_0000;
W1024R[500+180] = 16'b0000_0001_0000_0000;
W1024R[500+181] = 16'b0000_0001_0000_0000;
W1024R[500+182] = 16'b0000_0001_0000_0000;
W1024R[500+183] = 16'b0000_0001_0000_0000;
W1024R[500+184] = 16'b0000_0001_0000_0000;
W1024R[500+185] = 16'b0000_0001_0000_0000;
W1024R[500+186] = 16'b0000_0001_0000_0000;
W1024R[500+187] = 16'b0000_0001_0000_0000;
W1024R[500+188] = 16'b0000_0001_0000_0000;
W1024R[500+189] = 16'b0000_0001_0000_0000;
W1024R[500+190] = 16'b0000_0001_0000_0000;
W1024R[500+191] = 16'b0000_0001_0000_0000;
W1024R[500+192] = 16'b0000_0001_0000_0000;
W1024R[500+193] = 16'b0000_0001_0000_0000;
W1024R[500+194] = 16'b0000_0001_0000_0000;
W1024R[500+195] = 16'b0000_0001_0000_0000;
W1024R[500+196] = 16'b0000_0001_0000_0000;
W1024R[500+197] = 16'b0000_0001_0000_0000;
W1024R[500+198] = 16'b0000_0001_0000_0000;
W1024R[500+199] = 16'b0000_0001_0000_0000;

W1024R[600+100] = 16'b0000_0001_0000_0000;
W1024R[600+101] = 16'b0000_0001_0000_0000;
W1024R[600+102] = 16'b0000_0001_0000_0000;
W1024R[600+103] = 16'b0000_0001_0000_0000;
W1024R[600+104] = 16'b0000_0001_0000_0000;
W1024R[600+105] = 16'b0000_0001_0000_0000;
W1024R[600+106] = 16'b0000_0001_0000_0000;
W1024R[600+107] = 16'b0000_0001_0000_0000;
W1024R[600+108] = 16'b0000_0001_0000_0000;
W1024R[600+109] = 16'b0000_0001_0000_0000;
W1024R[600+110] = 16'b0000_0001_0000_0000;
W1024R[600+111] = 16'b0000_0001_0000_0000;
W1024R[600+112] = 16'b0000_0001_0000_0000;
W1024R[600+113] = 16'b0000_0001_0000_0000;
W1024R[600+114] = 16'b0000_0001_0000_0000;
W1024R[600+115] = 16'b0000_0001_0000_0000;
W1024R[600+116] = 16'b0000_0001_0000_0000;
W1024R[600+117] = 16'b0000_0001_0000_0000;
W1024R[600+118] = 16'b0000_0001_0000_0000;
W1024R[600+119] = 16'b0000_0001_0000_0000;
W1024R[600+120] = 16'b0000_0001_0000_0000;
W1024R[600+121] = 16'b0000_0001_0000_0000;
W1024R[600+122] = 16'b0000_0001_0000_0000;
W1024R[600+123] = 16'b0000_0001_0000_0000;
W1024R[600+124] = 16'b0000_0001_0000_0000;
W1024R[600+125] = 16'b0000_0001_0000_0000;
W1024R[600+126] = 16'b0000_0001_0000_0000;
W1024R[600+127] = 16'b0000_0001_0000_0000;
W1024R[600+128] = 16'b0000_0001_0000_0000;
W1024R[600+129] = 16'b0000_0001_0000_0000;
W1024R[600+130] = 16'b0000_0001_0000_0000;
W1024R[600+131] = 16'b0000_0001_0000_0000;
W1024R[600+132] = 16'b0000_0001_0000_0000;
W1024R[600+133] = 16'b0000_0001_0000_0000;
W1024R[600+134] = 16'b0000_0001_0000_0000;
W1024R[600+135] = 16'b0000_0001_0000_0000;
W1024R[600+136] = 16'b0000_0001_0000_0000;
W1024R[600+137] = 16'b0000_0001_0000_0000;
W1024R[600+138] = 16'b0000_0001_0000_0000;
W1024R[600+139] = 16'b0000_0001_0000_0000;
W1024R[600+140] = 16'b0000_0001_0000_0000;
W1024R[600+141] = 16'b0000_0001_0000_0000;
W1024R[600+142] = 16'b0000_0001_0000_0000;
W1024R[600+143] = 16'b0000_0001_0000_0000;
W1024R[600+144] = 16'b0000_0001_0000_0000;
W1024R[600+145] = 16'b0000_0001_0000_0000;
W1024R[600+146] = 16'b0000_0001_0000_0000;
W1024R[600+147] = 16'b0000_0001_0000_0000;
W1024R[600+148] = 16'b0000_0001_0000_0000;
W1024R[600+149] = 16'b0000_0001_0000_0000;
W1024R[600+150] = 16'b0000_0001_0000_0000;
W1024R[600+151] = 16'b0000_0001_0000_0000;
W1024R[600+152] = 16'b0000_0001_0000_0000;
W1024R[600+153] = 16'b0000_0001_0000_0000;
W1024R[600+154] = 16'b0000_0001_0000_0000;
W1024R[600+155] = 16'b0000_0001_0000_0000;
W1024R[600+156] = 16'b0000_0001_0000_0000;
W1024R[600+157] = 16'b0000_0001_0000_0000;
W1024R[600+158] = 16'b0000_0001_0000_0000;
W1024R[600+159] = 16'b0000_0001_0000_0000;
W1024R[600+160] = 16'b0000_0001_0000_0000;
W1024R[600+161] = 16'b0000_0001_0000_0000;
W1024R[600+162] = 16'b0000_0001_0000_0000;
W1024R[600+163] = 16'b0000_0001_0000_0000;
W1024R[600+164] = 16'b0000_0001_0000_0000;
W1024R[600+165] = 16'b0000_0001_0000_0000;
W1024R[600+166] = 16'b0000_0001_0000_0000;
W1024R[600+167] = 16'b0000_0001_0000_0000;
W1024R[600+168] = 16'b0000_0001_0000_0000;
W1024R[600+169] = 16'b0000_0001_0000_0000;
W1024R[600+170] = 16'b0000_0001_0000_0000;
W1024R[600+171] = 16'b0000_0001_0000_0000;
W1024R[600+172] = 16'b0000_0001_0000_0000;
W1024R[600+173] = 16'b0000_0001_0000_0000;
W1024R[600+174] = 16'b0000_0001_0000_0000;
W1024R[600+175] = 16'b0000_0001_0000_0000;
W1024R[600+176] = 16'b0000_0001_0000_0000;
W1024R[600+177] = 16'b0000_0001_0000_0000;
W1024R[600+178] = 16'b0000_0001_0000_0000;
W1024R[600+179] = 16'b0000_0001_0000_0000;
W1024R[600+180] = 16'b0000_0001_0000_0000;
W1024R[600+181] = 16'b0000_0001_0000_0000;
W1024R[600+182] = 16'b0000_0001_0000_0000;
W1024R[600+183] = 16'b0000_0001_0000_0000;
W1024R[600+184] = 16'b0000_0001_0000_0000;
W1024R[600+185] = 16'b0000_0001_0000_0000;
W1024R[600+186] = 16'b0000_0001_0000_0000;
W1024R[600+187] = 16'b0000_0001_0000_0000;
W1024R[600+188] = 16'b0000_0001_0000_0000;
W1024R[600+189] = 16'b0000_0001_0000_0000;
W1024R[600+190] = 16'b0000_0001_0000_0000;
W1024R[600+191] = 16'b0000_0001_0000_0000;
W1024R[600+192] = 16'b0000_0001_0000_0000;
W1024R[600+193] = 16'b0000_0001_0000_0000;
W1024R[600+194] = 16'b0000_0001_0000_0000;
W1024R[600+195] = 16'b0000_0001_0000_0000;
W1024R[600+196] = 16'b0000_0001_0000_0000;
W1024R[600+197] = 16'b0000_0001_0000_0000;
W1024R[600+198] = 16'b0000_0001_0000_0000;
W1024R[600+199] = 16'b0000_0001_0000_0000;

W1024R[700+100] = 16'b0000_0001_0000_0000;
W1024R[700+101] = 16'b0000_0001_0000_0000;
W1024R[700+102] = 16'b0000_0001_0000_0000;
W1024R[700+103] = 16'b0000_0001_0000_0000;
W1024R[700+104] = 16'b0000_0001_0000_0000;
W1024R[700+105] = 16'b0000_0001_0000_0000;
W1024R[700+106] = 16'b0000_0001_0000_0000;
W1024R[700+107] = 16'b0000_0001_0000_0000;
W1024R[700+108] = 16'b0000_0001_0000_0000;
W1024R[700+109] = 16'b0000_0001_0000_0000;
W1024R[700+110] = 16'b0000_0001_0000_0000;
W1024R[700+111] = 16'b0000_0001_0000_0000;
W1024R[700+112] = 16'b0000_0001_0000_0000;
W1024R[700+113] = 16'b0000_0001_0000_0000;
W1024R[700+114] = 16'b0000_0001_0000_0000;
W1024R[700+115] = 16'b0000_0001_0000_0000;
W1024R[700+116] = 16'b0000_0001_0000_0000;
W1024R[700+117] = 16'b0000_0001_0000_0000;
W1024R[700+118] = 16'b0000_0001_0000_0000;
W1024R[700+119] = 16'b0000_0001_0000_0000;
W1024R[700+120] = 16'b0000_0001_0000_0000;
W1024R[700+121] = 16'b0000_0001_0000_0000;
W1024R[700+122] = 16'b0000_0001_0000_0000;
W1024R[700+123] = 16'b0000_0001_0000_0000;
W1024R[700+124] = 16'b0000_0001_0000_0000;
W1024R[700+125] = 16'b0000_0001_0000_0000;
W1024R[700+126] = 16'b0000_0001_0000_0000;
W1024R[700+127] = 16'b0000_0001_0000_0000;
W1024R[700+128] = 16'b0000_0001_0000_0000;
W1024R[700+129] = 16'b0000_0001_0000_0000;
W1024R[700+130] = 16'b0000_0001_0000_0000;
W1024R[700+131] = 16'b0000_0001_0000_0000;
W1024R[700+132] = 16'b0000_0001_0000_0000;
W1024R[700+133] = 16'b0000_0001_0000_0000;
W1024R[700+134] = 16'b0000_0001_0000_0000;
W1024R[700+135] = 16'b0000_0001_0000_0000;
W1024R[700+136] = 16'b0000_0001_0000_0000;
W1024R[700+137] = 16'b0000_0001_0000_0000;
W1024R[700+138] = 16'b0000_0001_0000_0000;
W1024R[700+139] = 16'b0000_0001_0000_0000;
W1024R[700+140] = 16'b0000_0001_0000_0000;
W1024R[700+141] = 16'b0000_0001_0000_0000;
W1024R[700+142] = 16'b0000_0001_0000_0000;
W1024R[700+143] = 16'b0000_0001_0000_0000;
W1024R[700+144] = 16'b0000_0001_0000_0000;
W1024R[700+145] = 16'b0000_0001_0000_0000;
W1024R[700+146] = 16'b0000_0001_0000_0000;
W1024R[700+147] = 16'b0000_0001_0000_0000;
W1024R[700+148] = 16'b0000_0001_0000_0000;
W1024R[700+149] = 16'b0000_0001_0000_0000;
W1024R[700+150] = 16'b0000_0001_0000_0000;
W1024R[700+151] = 16'b0000_0001_0000_0000;
W1024R[700+152] = 16'b0000_0001_0000_0000;
W1024R[700+153] = 16'b0000_0001_0000_0000;
W1024R[700+154] = 16'b0000_0001_0000_0000;
W1024R[700+155] = 16'b0000_0001_0000_0000;
W1024R[700+156] = 16'b0000_0001_0000_0000;
W1024R[700+157] = 16'b0000_0001_0000_0000;
W1024R[700+158] = 16'b0000_0001_0000_0000;
W1024R[700+159] = 16'b0000_0001_0000_0000;
W1024R[700+160] = 16'b0000_0001_0000_0000;
W1024R[700+161] = 16'b0000_0001_0000_0000;
W1024R[700+162] = 16'b0000_0001_0000_0000;
W1024R[700+163] = 16'b0000_0001_0000_0000;
W1024R[700+164] = 16'b0000_0001_0000_0000;
W1024R[700+165] = 16'b0000_0001_0000_0000;
W1024R[700+166] = 16'b0000_0001_0000_0000;
W1024R[700+167] = 16'b0000_0001_0000_0000;
W1024R[700+168] = 16'b0000_0001_0000_0000;
W1024R[700+169] = 16'b0000_0001_0000_0000;
W1024R[700+170] = 16'b0000_0001_0000_0000;
W1024R[700+171] = 16'b0000_0001_0000_0000;
W1024R[700+172] = 16'b0000_0001_0000_0000;
W1024R[700+173] = 16'b0000_0001_0000_0000;
W1024R[700+174] = 16'b0000_0001_0000_0000;
W1024R[700+175] = 16'b0000_0001_0000_0000;
W1024R[700+176] = 16'b0000_0001_0000_0000;
W1024R[700+177] = 16'b0000_0001_0000_0000;
W1024R[700+178] = 16'b0000_0001_0000_0000;
W1024R[700+179] = 16'b0000_0001_0000_0000;
W1024R[700+180] = 16'b0000_0001_0000_0000;
W1024R[700+181] = 16'b0000_0001_0000_0000;
W1024R[700+182] = 16'b0000_0001_0000_0000;
W1024R[700+183] = 16'b0000_0001_0000_0000;
W1024R[700+184] = 16'b0000_0001_0000_0000;
W1024R[700+185] = 16'b0000_0001_0000_0000;
W1024R[700+186] = 16'b0000_0001_0000_0000;
W1024R[700+187] = 16'b0000_0001_0000_0000;
W1024R[700+188] = 16'b0000_0001_0000_0000;
W1024R[700+189] = 16'b0000_0001_0000_0000;
W1024R[700+190] = 16'b0000_0001_0000_0000;
W1024R[700+191] = 16'b0000_0001_0000_0000;
W1024R[700+192] = 16'b0000_0001_0000_0000;
W1024R[700+193] = 16'b0000_0001_0000_0000;
W1024R[700+194] = 16'b0000_0001_0000_0000;
W1024R[700+195] = 16'b0000_0001_0000_0000;
W1024R[700+196] = 16'b0000_0001_0000_0000;
W1024R[700+197] = 16'b0000_0001_0000_0000;
W1024R[700+198] = 16'b0000_0001_0000_0000;
W1024R[700+199] = 16'b0000_0001_0000_0000;

W1024R[800+100] = 16'b0000_0001_0000_0000;
W1024R[800+101] = 16'b0000_0001_0000_0000;
W1024R[800+102] = 16'b0000_0001_0000_0000;
W1024R[800+103] = 16'b0000_0001_0000_0000;
W1024R[800+104] = 16'b0000_0001_0000_0000;
W1024R[800+105] = 16'b0000_0001_0000_0000;
W1024R[800+106] = 16'b0000_0001_0000_0000;
W1024R[800+107] = 16'b0000_0001_0000_0000;
W1024R[800+108] = 16'b0000_0001_0000_0000;
W1024R[800+109] = 16'b0000_0001_0000_0000;
W1024R[800+110] = 16'b0000_0001_0000_0000;
W1024R[800+111] = 16'b0000_0001_0000_0000;
W1024R[800+112] = 16'b0000_0001_0000_0000;
W1024R[800+113] = 16'b0000_0001_0000_0000;
W1024R[800+114] = 16'b0000_0001_0000_0000;
W1024R[800+115] = 16'b0000_0001_0000_0000;
W1024R[800+116] = 16'b0000_0001_0000_0000;
W1024R[800+117] = 16'b0000_0001_0000_0000;
W1024R[800+118] = 16'b0000_0001_0000_0000;
W1024R[800+119] = 16'b0000_0001_0000_0000;
W1024R[800+120] = 16'b0000_0001_0000_0000;
W1024R[800+121] = 16'b0000_0001_0000_0000;
W1024R[800+122] = 16'b0000_0001_0000_0000;
W1024R[800+123] = 16'b0000_0001_0000_0000;
W1024R[800+124] = 16'b0000_0001_0000_0000;
W1024R[800+125] = 16'b0000_0001_0000_0000;
W1024R[800+126] = 16'b0000_0001_0000_0000;
W1024R[800+127] = 16'b0000_0001_0000_0000;
W1024R[800+128] = 16'b0000_0001_0000_0000;
W1024R[800+129] = 16'b0000_0001_0000_0000;
W1024R[800+130] = 16'b0000_0001_0000_0000;
W1024R[800+131] = 16'b0000_0001_0000_0000;
W1024R[800+132] = 16'b0000_0001_0000_0000;
W1024R[800+133] = 16'b0000_0001_0000_0000;
W1024R[800+134] = 16'b0000_0001_0000_0000;
W1024R[800+135] = 16'b0000_0001_0000_0000;
W1024R[800+136] = 16'b0000_0001_0000_0000;
W1024R[800+137] = 16'b0000_0001_0000_0000;
W1024R[800+138] = 16'b0000_0001_0000_0000;
W1024R[800+139] = 16'b0000_0001_0000_0000;
W1024R[800+140] = 16'b0000_0001_0000_0000;
W1024R[800+141] = 16'b0000_0001_0000_0000;
W1024R[800+142] = 16'b0000_0001_0000_0000;
W1024R[800+143] = 16'b0000_0001_0000_0000;
W1024R[800+144] = 16'b0000_0001_0000_0000;
W1024R[800+145] = 16'b0000_0001_0000_0000;
W1024R[800+146] = 16'b0000_0001_0000_0000;
W1024R[800+147] = 16'b0000_0001_0000_0000;
W1024R[800+148] = 16'b0000_0001_0000_0000;
W1024R[800+149] = 16'b0000_0001_0000_0000;
W1024R[800+150] = 16'b0000_0001_0000_0000;
W1024R[800+151] = 16'b0000_0001_0000_0000;
W1024R[800+152] = 16'b0000_0001_0000_0000;
W1024R[800+153] = 16'b0000_0001_0000_0000;
W1024R[800+154] = 16'b0000_0001_0000_0000;
W1024R[800+155] = 16'b0000_0001_0000_0000;
W1024R[800+156] = 16'b0000_0001_0000_0000;
W1024R[800+157] = 16'b0000_0001_0000_0000;
W1024R[800+158] = 16'b0000_0001_0000_0000;
W1024R[800+159] = 16'b0000_0001_0000_0000;
W1024R[800+160] = 16'b0000_0001_0000_0000;
W1024R[800+161] = 16'b0000_0001_0000_0000;
W1024R[800+162] = 16'b0000_0001_0000_0000;
W1024R[800+163] = 16'b0000_0001_0000_0000;
W1024R[800+164] = 16'b0000_0001_0000_0000;
W1024R[800+165] = 16'b0000_0001_0000_0000;
W1024R[800+166] = 16'b0000_0001_0000_0000;
W1024R[800+167] = 16'b0000_0001_0000_0000;
W1024R[800+168] = 16'b0000_0001_0000_0000;
W1024R[800+169] = 16'b0000_0001_0000_0000;
W1024R[800+170] = 16'b0000_0001_0000_0000;
W1024R[800+171] = 16'b0000_0001_0000_0000;
W1024R[800+172] = 16'b0000_0001_0000_0000;
W1024R[800+173] = 16'b0000_0001_0000_0000;
W1024R[800+174] = 16'b0000_0001_0000_0000;
W1024R[800+175] = 16'b0000_0001_0000_0000;
W1024R[800+176] = 16'b0000_0001_0000_0000;
W1024R[800+177] = 16'b0000_0001_0000_0000;
W1024R[800+178] = 16'b0000_0001_0000_0000;
W1024R[800+179] = 16'b0000_0001_0000_0000;
W1024R[800+180] = 16'b0000_0001_0000_0000;
W1024R[800+181] = 16'b0000_0001_0000_0000;
W1024R[800+182] = 16'b0000_0001_0000_0000;
W1024R[800+183] = 16'b0000_0001_0000_0000;
W1024R[800+184] = 16'b0000_0001_0000_0000;
W1024R[800+185] = 16'b0000_0001_0000_0000;
W1024R[800+186] = 16'b0000_0001_0000_0000;
W1024R[800+187] = 16'b0000_0001_0000_0000;
W1024R[800+188] = 16'b0000_0001_0000_0000;
W1024R[800+189] = 16'b0000_0001_0000_0000;
W1024R[800+190] = 16'b0000_0001_0000_0000;
W1024R[800+191] = 16'b0000_0001_0000_0000;
W1024R[800+192] = 16'b0000_0001_0000_0000;
W1024R[800+193] = 16'b0000_0001_0000_0000;
W1024R[800+194] = 16'b0000_0001_0000_0000;
W1024R[800+195] = 16'b0000_0001_0000_0000;
W1024R[800+196] = 16'b0000_0001_0000_0000;
W1024R[800+197] = 16'b0000_0001_0000_0000;
W1024R[800+198] = 16'b0000_0001_0000_0000;
W1024R[800+199] = 16'b0000_0001_0000_0000;

W1024R[1000] = 16'b0000_0001_0000_0000;
W1024R[1001] = 16'b0000_0001_0000_0000;
W1024R[1002] = 16'b0000_0001_0000_0000;
W1024R[1003] = 16'b0000_0001_0000_0000;
W1024R[1004] = 16'b0000_0001_0000_0000;
W1024R[1005] = 16'b0000_0001_0000_0000;
W1024R[1006] = 16'b0000_0001_0000_0000;
W1024R[1007] = 16'b0000_0001_0000_0000;
W1024R[1008] = 16'b0000_0001_0000_0000;
W1024R[1009] = 16'b0000_0001_0000_0000;
W1024R[1010] = 16'b0000_0001_0000_0000;
W1024R[1011] = 16'b0000_0001_0000_0000;
W1024R[1012] = 16'b0000_0001_0000_0000;
W1024R[1013] = 16'b0000_0001_0000_0000;
W1024R[1014] = 16'b0000_0001_0000_0000;
W1024R[1015] = 16'b0000_0001_0000_0000;
W1024R[1016] = 16'b0000_0001_0000_0000;
W1024R[1017] = 16'b0000_0001_0000_0000;
W1024R[1018] = 16'b0000_0001_0000_0000;
W1024R[1019] = 16'b0000_0001_0000_0000;
W1024R[1020] = 16'b0000_0001_0000_0000;
W1024R[1021] = 16'b0000_0001_0000_0000;
W1024R[1022] = 16'b0000_0001_0000_0000;
W1024R[1023] = 16'b0000_0001_0000_0000;
            
            //其他1023个点交给你喽@李孟锡
        end    //rstn
        else begin
             case(current_state)
             S0:begin
                if(req_input_c == 1'b1) next_state = S1;    //从复位态到输入态的方法
                else next_state = S0;
                ans_input2 = 1'b0;
                en_input = 1'b0;
                req_output = 1'b0;    //控制信号
                en_output = 1'b0;
                input_count = 10'b00000_00000;    //为输入级做初始化
                end    //S0
             S1:begin
                req_output = 1'b0;    //控制信号
                en_output = 1'b0;
                if(req_input_c == 1'b1) begin
                    en_input = 1'b1;
                    ans_input2 = 1'b1;
                end
                if(input_count == 10'b11111_11111) next_state = S2;    //输入态-->处理态
                else next_state = S1;
                ji = 4'b0000;
                position = 10'b00000_00000;    //为运算级做初始化
                end    //S1
             
             S2:begin
                ans_input2 = 1'b0;
                en_input = 1'b0;
                req_output = 1'b0;    //控制信号
                en_output = 1'b0;
                output_count = 10'b00000_00000;
                if(ji == 4'b0000) begin
                    next_ji = 4'b0001;
                    next_position = 10'b00000_00000;
                    next_state = S2;
                end
                if(position < 10'b11111_11111) begin
                next_ji = ji;
                next_position = position + 10'b00000_00001;
                next_state = S2;
                end
                else begin
                    if(ji < 4'b1010) begin
                         next_position = 10'b00000_00000;
                         next_ji = ji + 4'b0001;
                         next_state = S2;
                    end
                    else begin
                        next_position = 10'b00000_00000;
                        next_ji = 4'b0000;
                        next_state = S3;    //ji=10,position计满，进入下个状态
                    end
                end    //else
                case(ji)
                4'b0000:begin    //第零级,只有一个周期，为了为第一级做缓冲
                e <= fft0R[0];    //在当前位置要考虑下一位置的运算
                f <= fft0J[0];
                a <= fft0R[1];
                b <= fft0J[1];
                c <= W1024R[0];
                d <= W1024J[0];
                end    //0000
                4'b0001:begin
                if(position == 10'b11111_11111) begin
                    e <= fft1R[0];    //最后一个position为下一级缓冲
                    f <= fft1J[0];
                    a <= fft1R[2];
                    b <= fft1J[2];
                    c <= W1024R[0];
                    d <= W1024J[0];
                end    //if
                else begin
                    if(position[0] == 1'b0) begin
                        e <= fft0R[position_plus];    //常规操作：同址运算
                        f <= fft0J[position_plus];    //position+1为同址
                        a <= fft0R[position_plus+1];    //position+1+N/2为蝶形运算另一个操作数
                        b <= fft0J[position_plus+1];
                        c <= W1024R[position_plus[0]*512];    //旋转因子相对确定
                        d <= W1024J[position_plus[0]*512];
                    end
                    else begin
                        e <= fft0R[position_plus-1];    //非常规操作：同址旋转+
                        f <= fft0J[position_plus-1];
                        a <= fft0R[position_plus];
                        b <= fft0J[position_plus];
                        c <= W1024R[position_plus[0]*512];
                        d <= W1024J[position_plus[0]*512];
                    end
                end    //else
                end    //0001
                4'b0010:begin
                if(position == 10'b11111_11111) begin
                    e <= fft2R[0];    //最后一个position为下一级缓冲
                    f <= fft2J[0];
                    a <= fft2R[4];
                    b <= fft2J[4];
                    c <= W1024R[0];
                    d <= W1024J[0];
                end    //if
                else begin
                    if(position[1] == 1'b0) begin
                        e <= fft1R[position_plus];
                        f <= fft1J[position_plus];
                        a <= fft1R[position_plus+2];
                        b <= fft1J[position_plus+2];
                        c <= W1024R[position_plus[1:0]*256];
                        d <= W1024J[position_plus[1:0]*256];
                    end
                    else begin
                        e <= fft1R[position_plus-2];
                        f <= fft1J[position_plus-2];
                        a <= fft1R[position_plus];
                        b <= fft1J[position_plus];
                        c <= W1024R[position_plus[1:0]*256];
                        d <= W1024J[position_plus[1:0]*256];
                    end
                end    //else
                end
                4'b0011:begin
                if(position == 10'b11111_11111) begin
                    e <= fft3R[0];    //最后一个position为下一级缓冲
                    f <= fft3J[0];
                    a <= fft3R[8];
                    b <= fft3J[8];
                    c <= W1024R[0];
                    d <= W1024J[0];
                end    //if
                else begin
                    if(position[2] == 1'b0) begin
                        e <= fft2R[position_plus];
                        f <= fft2J[position_plus];
                        a <= fft2R[position_plus+4];
                        b <= fft2J[position_plus+4];
                        c <= W1024R[position_plus[2:0]*128];
                        d <= W1024J[position_plus[2:0]*128];
                    end
                    else begin
                        e <= fft2R[position_plus-4];
                        f <= fft2J[position_plus-4];
                        a <= fft2R[position_plus];
                        b <= fft2J[position_plus];
                        c <= W1024R[position_plus[2:0]*128];
                        d <= W1024J[position_plus[2:0]*128];
                    end
                end    //else
                end
                4'b0100:begin
                if(position == 10'b11111_11111) begin
                    e <= fft4R[0];    //最后一个position为下一级缓冲
                    f <= fft4J[0];
                    a <= fft4R[16];
                    b <= fft4J[16];
                    c <= W1024R[0];
                    d <= W1024J[0];
                end    //if
                else begin
                    if(position[3] == 1'b0) begin
                        e <= fft3R[position_plus];
                        f <= fft3J[position_plus];
                        a <= fft3R[position_plus+8];
                        b <= fft3J[position_plus+8];
                        c <= W1024R[position_plus[3:0]*64];
                        d <= W1024J[position_plus[3:0]*64];
                    end
                    else begin
                        e <= fft3R[position_plus-8];
                        f <= fft3J[position_plus-8];
                        a <= fft3R[position_plus];
                        b <= fft3J[position_plus];
                        c <= W1024R[position_plus[3:0]*64];
                        d <= W1024J[position_plus[3:0]*64];
                    end
                end    //else
                end
                4'b0101:begin
                if(position == 10'b11111_11111) begin
                    e <= fft5R[0];    //最后一个position为下一级缓冲
                    f <= fft5J[0];
                    a <= fft5R[32];
                    b <= fft5J[32];
                    c <= W1024R[0];
                    d <= W1024J[0];
                end    //if
                else begin
                    if(position[4] == 1'b0) begin
                        e <= fft4R[position_plus];
                        f <= fft4J[position_plus];
                        a <= fft4R[position_plus+16];
                        b <= fft4J[position_plus+16];
                        c <= W1024R[position_plus[4:0]*32];
                        d <= W1024J[position_plus[4:0]*32];
                    end
                    else begin
                        e <= fft4R[position_plus-16];
                        f <= fft4J[position_plus-16];
                        a <= fft4R[position_plus];
                        b <= fft4J[position_plus];
                        c <= W1024R[position_plus[4:0]*32];
                        d <= W1024J[position_plus[4:0]*32];
                    end
                end    //else
                end
                4'b0110:begin
                if(position == 10'b11111_11111) begin
                    e <= fft6R[0];    //最后一个position为下一级缓冲
                    f <= fft6J[0];
                    a <= fft6R[64];
                    b <= fft6J[64];
                    c <= W1024R[0];
                    d <= W1024J[0];
                end    //if
                else begin
                    if(position[5] == 1'b0) begin
                        e <= fft5R[position_plus];
                        f <= fft5J[position_plus];
                        a <= fft5R[position_plus+32];
                        b <= fft5J[position_plus+32];
                        c <= W1024R[position_plus[5:0]*16];
                        d <= W1024J[position_plus[5:0]*16];
                    end
                    else begin
                        e <= fft5R[position_plus-32];
                        f <= fft5J[position_plus-32];
                        a <= fft5R[position_plus];
                        b <= fft5J[position_plus];
                        c <= W1024R[position_plus[5:0]*16];
                        d <= W1024J[position_plus[5:0]*16];
                    end
                end    //else
                end
                4'b0111:begin
                if(position == 10'b11111_11111) begin
                    e <= fft7R[0];    //最后一个position为下一级缓冲
                    f <= fft7J[0];
                    a <= fft7R[128];
                    b <= fft7J[128];
                    c <= W1024R[0];
                    d <= W1024J[0];
                end    //if
                else begin
                    if(position[6] == 1'b0) begin
                        e <= fft6R[position_plus];
                        f <= fft6J[position_plus];
                        a <= fft6R[position_plus+64];
                        b <= fft6J[position_plus+64];
                        c <= W1024R[position_plus[6:0]*8];
                        d <= W1024J[position_plus[6:0]*8];
                    end
                    else begin
                        e <= fft6R[position_plus-64];
                        f <= fft6J[position_plus-64];
                        a <= fft6R[position_plus];
                        b <= fft6J[position_plus];
                        c <= W1024R[position_plus[6:0]*8];
                        d <= W1024J[position_plus[6:0]*8];
                    end
                end    //else
                end
                4'b1000:begin
                if(position == 10'b11111_11111) begin
                    e <= fft8R[0];    //最后一个position为下一级缓冲
                    f <= fft8J[0];
                    a <= fft8R[256];
                    b <= fft8J[256];
                    c <= W1024R[0];
                    d <= W1024J[0];
                end    //if
                else begin
                    if(position[7] == 1'b0) begin
                        e <= fft7R[position_plus];
                        f <= fft7J[position_plus];
                        a <= fft7R[position_plus+128];
                        b <= fft7J[position_plus+128];
                        c <= W1024R[position_plus[7:0]*4];
                        d <= W1024J[position_plus[7:0]*4];
                    end
                    else begin
                        e <= fft7R[position_plus-128];
                        f <= fft7J[position_plus-128];
                        a <= fft7R[position_plus];
                        b <= fft7J[position_plus];
                        c <= W1024R[position_plus[7:0]*4];
                        d <= W1024J[position_plus[7:0]*4];
                    end
                end    //else
                end
                4'b1001:begin
                if(position == 10'b11111_11111) begin
                    e <= fft9R[0];    //最后一个position为下一级缓冲
                    f <= fft9J[0];
                    a <= fft9R[512];
                    b <= fft9J[512];
                    c <= W1024R[0];
                    d <= W1024J[0];
                end    //if
                else begin
                    if(position[8] == 1'b0) begin
                        e <= fft8R[position_plus];
                        f <= fft8J[position_plus];
                        a <= fft8R[position_plus+256];
                        b <= fft8J[position_plus+256];
                        c <= W1024R[position_plus[8:0]*2];
                        d <= W1024J[position_plus[8:0]*2];
                    end
                    else begin
                        e <= fft8R[position_plus-256];
                        f <= fft8J[position_plus-256];
                        a <= fft8R[position_plus];
                        b <= fft8J[position_plus];
                        c <= W1024R[position_plus[8:0]*2];
                        d <= W1024J[position_plus[8:0]*2];
                    end
                end    //else
                end
                4'b1010:begin
                if(position[9] == 1'b0) begin
                    e <= fft9R[position_plus];
                    f <= fft9J[position_plus];
                    a <= fft9R[position_plus+512];
                    b <= fft9J[position_plus+512];
                    c <= W1024R[position_plus[9:0]];
                    d <= W1024J[position_plus[9:0]];
                end
                else begin
                    e <= fft8R[position_plus-512];
                    f <= fft8J[position_plus-512];
                    a <= fft8R[position_plus];
                    b <= fft8J[position_plus];
                    c <= W1024R[position_plus[9:0]];
                    d <= W1024J[position_plus[9:0]];
                end
                end
                default:begin
                
                end
                endcase
                end    //S2
             S3:begin
                en_input = 1'b0;
                ans_input2 = 1'b0;
                req_output = 1'b1;
                en_output = 1'b0;
                if(output_count == 10'b11111_11111) begin
                    next_state = S0;
                end
                end
             endcase
        end    //else
    end
    
    always @(*) begin    //组合逻辑将wire连到寄存器（暂时保留）
        data_oR = data_oR_c;
        data_oJ = data_oJ_c;
        req_o = req_o_c;
        ans_o = ans_input1_c;
        position_plus = position+1;
    end
    
fft_input fft_input
     (.rstn(rstn),    //.端口名（线网名）
      .req_i(req_i),    //请求输入（从外adc）
      .data_i(data_i),    //数据输入（从外adc）
      .ans_i(ans_input2),    //反馈（从FPGA）
      .en(en_input),    //使能（从FPGA）
      .req_o(req_input_c),    //请求（到FPGA）
      .ans_o(ans_input1_c),    //反馈告知外部
      .data_o(data_input_c)    //数据输出（到FPGA）
      );
      
fft_output fft_output
     (.rstn(rstn),
      .req_i(req_output),    //请求输入（从FPGA）
      .ans_i(ans_i),    //反馈输入（从MCU）
      .en(en_output),    //使能
      .data_iR(),    //数据输出（从FPGA）
      .data_iJ(),
      .req_o(req_o_c),    //请求输出（到MCU）
      .ans_o(ans_output1_c),    //反馈输出（到FPGA）
      .data_oR(data_oR_c),    //数据输出（到MCU）
      .data_oJ(data_oJ_c)
      );
MAC MAC
    (.rstn(rstn),
     .a(a),
     .b(b),
     .c(c),
     .d(d),
     .e(e),
     .f(f),
     .R(R),
     .J(J),
     .over_a(over_a),
     .over_m(over_m)
     );
endmodule
